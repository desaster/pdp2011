
--
-- Copyright (c) 2008-2020 Sytse van Slooten
--
-- Permission is hereby granted to any person obtaining a copy of these VHDL source files and
-- other language source files and associated documentation files ("the materials") to use
-- these materials solely for personal, non-commercial purposes.
-- You are also granted permission to make changes to the materials, on the condition that this
-- copyright notice is retained unchanged.
--
-- The materials are distributed in the hope that they will be useful, but WITHOUT ANY WARRANTY;
-- without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.
--

-- $Revision$

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity xubr is
   port(
      base_addr : in std_logic_vector(17 downto 0);

      bus_addr_match : out std_logic;
      bus_addr : in std_logic_vector(17 downto 0);
      bus_dati : out std_logic_vector(15 downto 0);
      bus_dato : in std_logic_vector(15 downto 0);
      bus_control_dati : in std_logic;
      bus_control_dato : in std_logic;
      bus_control_datob : in std_logic;

      reset : in std_logic;
      clk : in std_logic
   );
end xubr;

architecture implementation of xubr is

signal base_addr_match : std_logic;

subtype u is std_logic_vector(7 downto 0);
type mem_type is array(0 to 4095) of u;

-- code base at 0

signal meme : mem_type := mem_type'(
u'(x"77"),u'(x"fc"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"df"),u'(x"e0"),u'(x"fe"),u'(x"c6"),u'(x"00"),u'(x"37"),u'(x"62"),u'(x"df"),u'(x"36"),u'(x"40"),u'(x"df"),u'(x"e0"),u'(x"42"),u'(x"df"),u'(x"40"),u'(x"66"),
u'(x"f7"),u'(x"ac"),u'(x"f7"),u'(x"02"),u'(x"f7"),u'(x"70"),u'(x"48"),u'(x"6c"),u'(x"6f"),u'(x"20"),u'(x"6f"),u'(x"6c"),u'(x"3a"),u'(x"78"),u'(x"2d"),u'(x"70"),
u'(x"20"),u'(x"74"),u'(x"35"),u'(x"20"),u'(x"65"),u'(x"6e"),u'(x"20"),u'(x"69"),u'(x"72"),u'(x"63"),u'(x"64"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"b2"),u'(x"1f"),
u'(x"fe"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"c0"),u'(x"03"),u'(x"1f"),u'(x"4a"),u'(x"04"),u'(x"df"),u'(x"02"),u'(x"4a"),u'(x"00"),u'(x"37"),u'(x"f2"),u'(x"f7"),
u'(x"e6"),u'(x"09"),u'(x"f7"),u'(x"28"),u'(x"f7"),u'(x"3e"),u'(x"04"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"f2"),u'(x"37"),u'(x"6e"),u'(x"f7"),u'(x"e0"),u'(x"06"),
u'(x"10"),u'(x"08"),u'(x"10"),u'(x"f7"),u'(x"5e"),u'(x"5d"),u'(x"f7"),u'(x"ec"),u'(x"63"),u'(x"6e"),u'(x"6f"),u'(x"20"),u'(x"65"),u'(x"64"),u'(x"65"),u'(x"64"),
u'(x"65"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"46"),u'(x"f7"),u'(x"5c"),u'(x"f7"),u'(x"a0"),u'(x"0f"),u'(x"f7"),u'(x"9b"),u'(x"0c"),u'(x"f7"),u'(x"96"),u'(x"09"),
u'(x"f7"),u'(x"91"),u'(x"06"),u'(x"f7"),u'(x"8c"),u'(x"03"),u'(x"f7"),u'(x"87"),u'(x"1e"),u'(x"f7"),u'(x"a6"),u'(x"72"),u'(x"73"),u'(x"6f"),u'(x"69"),u'(x"67"),
u'(x"6c"),u'(x"61"),u'(x"0a"),u'(x"f7"),u'(x"68"),u'(x"70"),u'(x"f7"),u'(x"63"),u'(x"6b"),u'(x"f7"),u'(x"5e"),u'(x"62"),u'(x"f7"),u'(x"59"),u'(x"5d"),u'(x"f7"),
u'(x"54"),u'(x"54"),u'(x"f7"),u'(x"4f"),u'(x"4f"),u'(x"f7"),u'(x"10"),u'(x"f7"),u'(x"40"),u'(x"0f"),u'(x"f7"),u'(x"64"),u'(x"72"),u'(x"73"),u'(x"6f"),u'(x"69"),
u'(x"67"),u'(x"6d"),u'(x"64"),u'(x"62"),u'(x"74"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"ea"),u'(x"f7"),u'(x"46"),u'(x"63"),u'(x"69"),u'(x"20"),u'(x"65"),u'(x"65"),
u'(x"0d"),u'(x"00"),u'(x"8a"),u'(x"f7"),u'(x"52"),u'(x"c0"),u'(x"4a"),u'(x"c0"),u'(x"f0"),u'(x"c0"),u'(x"02"),u'(x"77"),u'(x"00"),u'(x"c0"),u'(x"02"),u'(x"02"),
u'(x"77"),u'(x"f6"),u'(x"c0"),u'(x"03"),u'(x"02"),u'(x"77"),u'(x"ec"),u'(x"f7"),u'(x"0a"),u'(x"70"),u'(x"73"),u'(x"31"),u'(x"76"),u'(x"6c"),u'(x"65"),u'(x"77"),
u'(x"6f"),u'(x"67"),u'(x"3a"),u'(x"00"),u'(x"f7"),u'(x"56"),u'(x"48"),u'(x"08"),u'(x"f7"),u'(x"e8"),u'(x"0d"),u'(x"00"),u'(x"77"),u'(x"be"),u'(x"c1"),u'(x"48"),
u'(x"c1"),u'(x"20"),u'(x"04"),u'(x"1f"),u'(x"48"),u'(x"77"),u'(x"32"),u'(x"c1"),u'(x"10"),u'(x"02"),u'(x"77"),u'(x"16"),u'(x"1f"),u'(x"48"),u'(x"c1"),u'(x"f0"),
u'(x"77"),u'(x"8a"),u'(x"c1"),u'(x"c1"),u'(x"b0"),u'(x"41"),u'(x"c9"),u'(x"87"),u'(x"f7"),u'(x"a8"),u'(x"70"),u'(x"73"),u'(x"30"),u'(x"6e"),u'(x"6f"),u'(x"20"),
u'(x"20"),u'(x"f7"),u'(x"fc"),u'(x"48"),u'(x"02"),u'(x"f7"),u'(x"8e"),u'(x"0d"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"7e"),u'(x"70"),
u'(x"73"),u'(x"30"),u'(x"6e"),u'(x"6f"),u'(x"78"),u'(x"20"),u'(x"f7"),u'(x"d2"),u'(x"48"),u'(x"02"),u'(x"f7"),u'(x"64"),u'(x"0d"),u'(x"00"),u'(x"df"),u'(x"00"),
u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"54"),u'(x"70"),u'(x"73"),u'(x"30"),u'(x"63"),u'(x"64"),u'(x"20"),u'(x"65"),u'(x"20"),u'(x"63"),u'(x"62"),u'(x"3a"),u'(x"00"),
u'(x"f7"),u'(x"9e"),u'(x"48"),u'(x"08"),u'(x"f7"),u'(x"30"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"4c"),u'(x"58"),u'(x"f7"),u'(x"4e"),u'(x"54"),u'(x"df"),u'(x"00"),
u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"14"),u'(x"70"),u'(x"73"),u'(x"30"),u'(x"63"),u'(x"64"),u'(x"20"),u'(x"65"),u'(x"20"),u'(x"6d"),u'(x"3a"),u'(x"00"),u'(x"f7"),
u'(x"60"),u'(x"48"),u'(x"08"),u'(x"f7"),u'(x"f2"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"4c"),u'(x"0a"),u'(x"f7"),u'(x"4e"),u'(x"06"),u'(x"f7"),u'(x"e8"),u'(x"00"),
u'(x"00"),u'(x"d2"),u'(x"08"),u'(x"f7"),u'(x"d2"),u'(x"70"),u'(x"62"),u'(x"20"),u'(x"63"),u'(x"64"),u'(x"20"),u'(x"20"),u'(x"f7"),u'(x"26"),u'(x"d2"),u'(x"08"),
u'(x"f7"),u'(x"b8"),u'(x"0d"),u'(x"00"),u'(x"c0"),u'(x"e6"),u'(x"c0"),u'(x"16"),u'(x"05"),u'(x"c0"),u'(x"c0"),u'(x"d0"),u'(x"00"),u'(x"c8"),u'(x"87"),u'(x"df"),
u'(x"00"),u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"92"),u'(x"70"),u'(x"73"),u'(x"30"),u'(x"53"),u'(x"41"),u'(x"54"),u'(x"3a"),u'(x"00"),u'(x"f7"),u'(x"e4"),u'(x"48"),
u'(x"08"),u'(x"f7"),u'(x"76"),u'(x"0d"),u'(x"00"),u'(x"df"),u'(x"03"),u'(x"4a"),u'(x"f7"),u'(x"34"),u'(x"12"),u'(x"f7"),u'(x"01"),u'(x"2c"),u'(x"f7"),u'(x"34"),
u'(x"54"),u'(x"f7"),u'(x"30"),u'(x"50"),u'(x"f7"),u'(x"34"),u'(x"40"),u'(x"f7"),u'(x"30"),u'(x"3c"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),u'(x"df"),u'(x"00"),
u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"18"),u'(x"f7"),u'(x"60"),u'(x"03"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"1c"),
u'(x"70"),u'(x"73"),u'(x"30"),u'(x"53"),u'(x"4f"),u'(x"20"),u'(x"20"),u'(x"f7"),u'(x"70"),u'(x"48"),u'(x"08"),u'(x"f7"),u'(x"02"),u'(x"0d"),u'(x"00"),u'(x"37"),
u'(x"c6"),u'(x"df"),u'(x"02"),u'(x"4a"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),u'(x"f0"),u'(x"44"),u'(x"84"),u'(x"fe"),u'(x"06"),u'(x"5c"),u'(x"1a"),u'(x"1a"),
u'(x"64"),u'(x"1a"),u'(x"1a"),u'(x"1a"),u'(x"1a"),u'(x"1a"),u'(x"1a"),u'(x"7c"),u'(x"00"),u'(x"1a"),u'(x"3c"),u'(x"f0"),u'(x"14"),u'(x"7a"),u'(x"e0"),u'(x"32"),
u'(x"62"),u'(x"d8"),u'(x"d4"),u'(x"f8"),u'(x"26"),u'(x"68"),u'(x"bc"),u'(x"ca"),u'(x"d8"),u'(x"02"),u'(x"2c"),u'(x"3a"),u'(x"48"),u'(x"56"),u'(x"64"),u'(x"72"),
u'(x"f7"),u'(x"98"),u'(x"66"),u'(x"30"),u'(x"2d"),u'(x"6e"),u'(x"6f"),u'(x"0d"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"7e"),u'(x"66"),
u'(x"31"),u'(x"2d"),u'(x"6c"),u'(x"61"),u'(x"20"),u'(x"6e"),u'(x"20"),u'(x"74"),u'(x"72"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"5c"),
u'(x"66"),u'(x"32"),u'(x"2d"),u'(x"72"),u'(x"61"),u'(x"20"),u'(x"65"),u'(x"61"),u'(x"6c"),u'(x"20"),u'(x"68"),u'(x"73"),u'(x"63"),u'(x"6c"),u'(x"61"),u'(x"64"),
u'(x"65"),u'(x"73"),u'(x"00"),u'(x"f7"),u'(x"64"),u'(x"f7"),u'(x"56"),u'(x"00"),u'(x"01"),u'(x"f7"),u'(x"26"),u'(x"3a"),u'(x"f7"),u'(x"48"),u'(x"01"),u'(x"01"),
u'(x"f7"),u'(x"18"),u'(x"3a"),u'(x"f7"),u'(x"3a"),u'(x"fe"),u'(x"01"),u'(x"f7"),u'(x"0a"),u'(x"3a"),u'(x"f7"),u'(x"2c"),u'(x"ff"),u'(x"01"),u'(x"f7"),u'(x"fc"),
u'(x"3a"),u'(x"f7"),u'(x"1e"),u'(x"fc"),u'(x"01"),u'(x"f7"),u'(x"ee"),u'(x"3a"),u'(x"f7"),u'(x"10"),u'(x"fd"),u'(x"01"),u'(x"f7"),u'(x"e0"),u'(x"0d"),u'(x"00"),
u'(x"f7"),u'(x"3c"),u'(x"0e"),u'(x"f7"),u'(x"37"),u'(x"09"),u'(x"f7"),u'(x"2e"),u'(x"04"),u'(x"f7"),u'(x"29"),u'(x"ff"),u'(x"f7"),u'(x"20"),u'(x"fa"),u'(x"f7"),
u'(x"1b"),u'(x"f5"),u'(x"f7"),u'(x"06"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"a8"),u'(x"66"),u'(x"33"),u'(x"2d"),u'(x"6e"),u'(x"20"),u'(x"70"),
u'(x"66"),u'(x"6e"),u'(x"74"),u'(x"6f"),u'(x"0d"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"84"),u'(x"66"),u'(x"34"),u'(x"2d"),u'(x"72"),
u'(x"61"),u'(x"20"),u'(x"68"),u'(x"73"),u'(x"63"),u'(x"6c"),u'(x"61"),u'(x"64"),u'(x"65"),u'(x"73"),u'(x"00"),u'(x"f7"),u'(x"94"),u'(x"f7"),u'(x"3a"),u'(x"94"),
u'(x"f7"),u'(x"35"),u'(x"8f"),u'(x"f7"),u'(x"30"),u'(x"8a"),u'(x"f7"),u'(x"2b"),u'(x"85"),u'(x"f7"),u'(x"26"),u'(x"80"),u'(x"f7"),u'(x"21"),u'(x"7b"),u'(x"f7"),
u'(x"62"),u'(x"d4"),u'(x"06"),u'(x"f7"),u'(x"32"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"7c"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"1e"),u'(x"66"),
u'(x"35"),u'(x"2d"),u'(x"77"),u'(x"69"),u'(x"65"),u'(x"70"),u'(x"79"),u'(x"69"),u'(x"61"),u'(x"20"),u'(x"64"),u'(x"72"),u'(x"73"),u'(x"20"),u'(x"f7"),u'(x"2e"),
u'(x"f7"),u'(x"30"),u'(x"d2"),u'(x"f7"),u'(x"2b"),u'(x"cd"),u'(x"f7"),u'(x"26"),u'(x"c8"),u'(x"f7"),u'(x"21"),u'(x"c3"),u'(x"f7"),u'(x"1c"),u'(x"be"),u'(x"f7"),
u'(x"17"),u'(x"b9"),u'(x"f7"),u'(x"fc"),u'(x"78"),u'(x"06"),u'(x"f7"),u'(x"cc"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"66"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),
u'(x"f7"),u'(x"b8"),u'(x"66"),u'(x"36"),u'(x"2d"),u'(x"72"),u'(x"61"),u'(x"20"),u'(x"75"),u'(x"74"),u'(x"63"),u'(x"73"),u'(x"20"),u'(x"64"),u'(x"72"),u'(x"73"),
u'(x"20"),u'(x"69"),u'(x"74"),u'(x"0a"),u'(x"f7"),u'(x"c2"),u'(x"c0"),u'(x"c7"),u'(x"c0"),u'(x"0a"),u'(x"0a"),u'(x"37"),u'(x"c0"),u'(x"c0"),u'(x"02"),u'(x"f7"),
u'(x"ca"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"66"),u'(x"66"),u'(x"37"),u'(x"2d"),u'(x"77"),u'(x"69"),
u'(x"65"),u'(x"6d"),u'(x"6c"),u'(x"69"),u'(x"61"),u'(x"74"),u'(x"61"),u'(x"64"),u'(x"65"),u'(x"73"),u'(x"6c"),u'(x"73"),u'(x"20"),u'(x"f7"),u'(x"70"),u'(x"c0"),
u'(x"75"),u'(x"37"),u'(x"76"),u'(x"c0"),u'(x"0c"),u'(x"f7"),u'(x"10"),u'(x"3a"),u'(x"20"),u'(x"00"),u'(x"00"),u'(x"f7"),u'(x"22"),u'(x"63"),u'(x"65"),u'(x"72"),
u'(x"64"),u'(x"c0"),u'(x"0a"),u'(x"69"),u'(x"f7"),u'(x"f2"),u'(x"36"),u'(x"20"),u'(x"00"),u'(x"00"),u'(x"f7"),u'(x"1e"),u'(x"f7"),u'(x"66"),u'(x"dc"),u'(x"02"),
u'(x"f7"),u'(x"f8"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"f0"),u'(x"66"),u'(x"37"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"f7"),u'(x"06"),u'(x"de"),
u'(x"0c"),u'(x"f7"),u'(x"d6"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"ce"),u'(x"66"),u'(x"37"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"f7"),u'(x"e4"),
u'(x"ea"),u'(x"0c"),u'(x"f7"),u'(x"b4"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"ac"),u'(x"66"),u'(x"37"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"f7"),
u'(x"c2"),u'(x"f6"),u'(x"0c"),u'(x"f7"),u'(x"92"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"8a"),u'(x"66"),u'(x"37"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"20"),
u'(x"f7"),u'(x"a0"),u'(x"02"),u'(x"0c"),u'(x"f7"),u'(x"70"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"68"),u'(x"66"),u'(x"37"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"20"),
u'(x"20"),u'(x"f7"),u'(x"7e"),u'(x"0e"),u'(x"0c"),u'(x"f7"),u'(x"4e"),u'(x"0d"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),u'(x"df"),u'(x"00"),u'(x"48"),
u'(x"87"),u'(x"f7"),u'(x"36"),u'(x"66"),u'(x"31"),u'(x"20"),u'(x"20"),u'(x"65"),u'(x"64"),u'(x"72"),u'(x"6e"),u'(x"20"),u'(x"6f"),u'(x"6d"),u'(x"74"),u'(x"0d"),
u'(x"00"),u'(x"f7"),u'(x"48"),u'(x"f7"),u'(x"ec"),u'(x"90"),u'(x"f7"),u'(x"e4"),u'(x"8c"),u'(x"f7"),u'(x"e2"),u'(x"87"),u'(x"f7"),u'(x"de"),u'(x"82"),u'(x"f7"),
u'(x"e0"),u'(x"7e"),u'(x"f7"),u'(x"d8"),u'(x"7a"),u'(x"f7"),u'(x"d6"),u'(x"75"),u'(x"f7"),u'(x"d2"),u'(x"70"),u'(x"f7"),u'(x"48"),u'(x"1c"),u'(x"0c"),u'(x"f7"),
u'(x"da"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"0c"),u'(x"4e"),u'(x"f7"),u'(x"5e"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"c0"),u'(x"66"),u'(x"31"),
u'(x"20"),u'(x"20"),u'(x"72"),u'(x"74"),u'(x"20"),u'(x"69"),u'(x"67"),u'(x"66"),u'(x"72"),u'(x"61"),u'(x"20"),u'(x"f7"),u'(x"d4"),u'(x"f7"),u'(x"0c"),u'(x"1a"),
u'(x"f7"),u'(x"0a"),u'(x"f7"),u'(x"fa"),u'(x"1c"),u'(x"0c"),u'(x"f7"),u'(x"8c"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"04"),u'(x"5c"),u'(x"f7"),u'(x"01"),u'(x"56"),
u'(x"f7"),u'(x"fa"),u'(x"4e"),u'(x"f7"),u'(x"fc"),u'(x"48"),u'(x"c0"),u'(x"ef"),u'(x"37"),u'(x"44"),u'(x"f7"),u'(x"e8"),u'(x"40"),u'(x"f7"),u'(x"e4"),u'(x"42"),
u'(x"f7"),u'(x"01"),u'(x"3c"),u'(x"f7"),u'(x"da"),u'(x"34"),u'(x"f7"),u'(x"fc"),u'(x"2e"),u'(x"c0"),u'(x"cf"),u'(x"37"),u'(x"2a"),u'(x"f7"),u'(x"c8"),u'(x"26"),
u'(x"df"),u'(x"00"),u'(x"48"),u'(x"f7"),u'(x"0a"),u'(x"2a"),u'(x"f7"),u'(x"06"),u'(x"26"),u'(x"f7"),u'(x"0a"),u'(x"16"),u'(x"f7"),u'(x"06"),u'(x"12"),u'(x"f7"),
u'(x"f2"),u'(x"f8"),u'(x"f7"),u'(x"ee"),u'(x"f4"),u'(x"c0"),u'(x"ec"),u'(x"c0"),u'(x"f7"),u'(x"e4"),u'(x"e8"),u'(x"77"),u'(x"e2"),u'(x"f7"),u'(x"da"),u'(x"de"),
u'(x"77"),u'(x"d8"),u'(x"c0"),u'(x"f4"),u'(x"f7"),u'(x"d4"),u'(x"da"),u'(x"f7"),u'(x"d0"),u'(x"d6"),u'(x"c0"),u'(x"ce"),u'(x"c0"),u'(x"f7"),u'(x"c6"),u'(x"ca"),
u'(x"77"),u'(x"c4"),u'(x"f7"),u'(x"bc"),u'(x"c0"),u'(x"77"),u'(x"ba"),u'(x"c0"),u'(x"f4"),u'(x"87"),u'(x"f7"),u'(x"c4"),u'(x"66"),u'(x"31"),u'(x"20"),u'(x"20"),
u'(x"65"),u'(x"64"),u'(x"63"),u'(x"75"),u'(x"74"),u'(x"72"),u'(x"0d"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"a0"),u'(x"66"),u'(x"31"),
u'(x"20"),u'(x"20"),u'(x"65"),u'(x"64"),u'(x"61"),u'(x"64"),u'(x"63"),u'(x"65"),u'(x"72"),u'(x"63"),u'(x"75"),u'(x"74"),u'(x"72"),u'(x"0d"),u'(x"00"),u'(x"df"),
u'(x"00"),u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"72"),u'(x"66"),u'(x"31"),u'(x"20"),u'(x"20"),u'(x"65"),u'(x"64"),u'(x"6d"),u'(x"64"),u'(x"20"),u'(x"69"),u'(x"73"),
u'(x"00"),u'(x"f7"),u'(x"bc"),u'(x"72"),u'(x"02"),u'(x"f7"),u'(x"4e"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"78"),u'(x"f7"),u'(x"18"),u'(x"78"),u'(x"f7"),u'(x"8e"),
u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"30"),u'(x"66"),u'(x"31"),u'(x"20"),u'(x"20"),u'(x"72"),u'(x"74"),u'(x"20"),u'(x"6f"),u'(x"65"),u'(x"62"),
u'(x"74"),u'(x"20"),u'(x"f7"),u'(x"7a"),u'(x"72"),u'(x"02"),u'(x"f7"),u'(x"0c"),u'(x"20"),u'(x"3e"),u'(x"00"),u'(x"f7"),u'(x"34"),u'(x"f7"),u'(x"36"),u'(x"d2"),
u'(x"f7"),u'(x"5e"),u'(x"72"),u'(x"02"),u'(x"f7"),u'(x"f0"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"88"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"dc"),
u'(x"66"),u'(x"31"),u'(x"0d"),u'(x"00"),u'(x"87"),u'(x"f7"),u'(x"ce"),u'(x"66"),u'(x"31"),u'(x"0d"),u'(x"00"),u'(x"87"),u'(x"f7"),u'(x"c0"),u'(x"66"),u'(x"32"),
u'(x"20"),u'(x"20"),u'(x"75"),u'(x"70"),u'(x"69"),u'(x"74"),u'(x"72"),u'(x"61"),u'(x"20"),u'(x"65"),u'(x"6f"),u'(x"79"),u'(x"0a"),u'(x"df"),u'(x"00"),u'(x"48"),
u'(x"87"),u'(x"f7"),u'(x"96"),u'(x"66"),u'(x"32"),u'(x"20"),u'(x"20"),u'(x"6f"),u'(x"64"),u'(x"69"),u'(x"74"),u'(x"72"),u'(x"61"),u'(x"20"),u'(x"65"),u'(x"6f"),
u'(x"79"),u'(x"0a"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"6c"),u'(x"66"),u'(x"32"),u'(x"0d"),u'(x"00"),u'(x"87"),u'(x"f7"),u'(x"5e"),u'(x"66"),
u'(x"32"),u'(x"0d"),u'(x"00"),u'(x"87"),u'(x"f7"),u'(x"50"),u'(x"66"),u'(x"32"),u'(x"0d"),u'(x"00"),u'(x"87"),u'(x"f7"),u'(x"42"),u'(x"66"),u'(x"32"),u'(x"0d"),
u'(x"00"),u'(x"87"),u'(x"f7"),u'(x"34"),u'(x"66"),u'(x"32"),u'(x"0d"),u'(x"00"),u'(x"87"),u'(x"f7"),u'(x"26"),u'(x"66"),u'(x"32"),u'(x"0d"),u'(x"00"),u'(x"87"),
u'(x"37"),u'(x"48"),u'(x"f7"),u'(x"10"),u'(x"05"),u'(x"f7"),u'(x"08"),u'(x"02"),u'(x"77"),u'(x"8c"),u'(x"26"),u'(x"f7"),u'(x"fe"),u'(x"04"),u'(x"f7"),u'(x"f6"),
u'(x"fc"),u'(x"37"),u'(x"e6"),u'(x"f7"),u'(x"90"),u'(x"f7"),u'(x"00"),u'(x"fe"),u'(x"01"),u'(x"35"),u'(x"f7"),u'(x"d4"),u'(x"01"),u'(x"0a"),u'(x"f7"),u'(x"00"),
u'(x"ec"),u'(x"01"),u'(x"13"),u'(x"f7"),u'(x"01"),u'(x"c0"),u'(x"f7"),u'(x"52"),u'(x"f7"),u'(x"00"),u'(x"d8"),u'(x"02"),u'(x"37"),u'(x"b0"),u'(x"f7"),u'(x"ac"),
u'(x"f7"),u'(x"00"),u'(x"c8"),u'(x"02"),u'(x"f7"),u'(x"5c"),u'(x"f7"),u'(x"98"),u'(x"f7"),u'(x"a8"),u'(x"aa"),u'(x"0b"),u'(x"f7"),u'(x"9e"),u'(x"a0"),u'(x"07"),
u'(x"f7"),u'(x"98"),u'(x"92"),u'(x"f7"),u'(x"90"),u'(x"8a"),u'(x"08"),u'(x"f7"),u'(x"8a"),u'(x"84"),u'(x"f7"),u'(x"82"),u'(x"7c"),u'(x"77"),u'(x"88"),u'(x"80"),
u'(x"87"),u'(x"f7"),u'(x"58"),u'(x"40"),u'(x"20"),u'(x"00"),u'(x"00"),u'(x"f7"),u'(x"4c"),u'(x"44"),u'(x"20"),u'(x"00"),u'(x"00"),u'(x"37"),u'(x"64"),u'(x"87"),
u'(x"22"),u'(x"00"),u'(x"22"),u'(x"00"),u'(x"f7"),u'(x"58"),u'(x"03"),u'(x"f7"),u'(x"00"),u'(x"5a"),u'(x"f7"),u'(x"4a"),u'(x"30"),u'(x"f7"),u'(x"20"),u'(x"88"),
u'(x"20"),u'(x"00"),u'(x"00"),u'(x"f7"),u'(x"14"),u'(x"1e"),u'(x"20"),u'(x"00"),u'(x"00"),u'(x"f7"),u'(x"08"),u'(x"16"),u'(x"10"),u'(x"18"),u'(x"10"),u'(x"f7"),
u'(x"02"),u'(x"94"),u'(x"f6"),u'(x"87"),u'(x"22"),u'(x"00"),u'(x"26"),u'(x"66"),u'(x"a6"),u'(x"e6"),u'(x"26"),u'(x"c3"),u'(x"10"),u'(x"c1"),u'(x"0e"),u'(x"c1"),
u'(x"01"),u'(x"c2"),u'(x"08"),u'(x"c2"),u'(x"fc"),u'(x"c0"),u'(x"c3"),u'(x"10"),u'(x"02"),u'(x"c0"),u'(x"10"),u'(x"04"),u'(x"c4"),u'(x"01"),u'(x"01"),u'(x"01"),
u'(x"84"),u'(x"5f"),u'(x"40"),u'(x"9f"),u'(x"42"),u'(x"df"),u'(x"62"),u'(x"44"),u'(x"df"),u'(x"00"),u'(x"47"),u'(x"1f"),u'(x"46"),u'(x"f7"),u'(x"c4"),u'(x"2f"),
u'(x"37"),u'(x"c0"),u'(x"f7"),u'(x"90"),u'(x"78"),u'(x"17"),u'(x"f7"),u'(x"89"),u'(x"71"),u'(x"13"),u'(x"f7"),u'(x"82"),u'(x"6a"),u'(x"0f"),u'(x"f7"),u'(x"7b"),
u'(x"63"),u'(x"0b"),u'(x"f7"),u'(x"74"),u'(x"5c"),u'(x"07"),u'(x"f7"),u'(x"6d"),u'(x"55"),u'(x"03"),u'(x"f7"),u'(x"01"),u'(x"8a"),u'(x"f7"),u'(x"5a"),u'(x"48"),
u'(x"f7"),u'(x"55"),u'(x"43"),u'(x"f7"),u'(x"50"),u'(x"3e"),u'(x"f7"),u'(x"4b"),u'(x"39"),u'(x"f7"),u'(x"46"),u'(x"34"),u'(x"f7"),u'(x"41"),u'(x"2f"),u'(x"37"),
u'(x"60"),u'(x"f7"),u'(x"c0"),u'(x"18"),u'(x"f7"),u'(x"2a"),u'(x"13"),u'(x"04"),u'(x"84"),u'(x"84"),u'(x"c4"),u'(x"c4"),u'(x"c4"),u'(x"37"),u'(x"06"),u'(x"f7"),
u'(x"1c"),u'(x"60"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"42"),u'(x"c3"),u'(x"10"),u'(x"04"),u'(x"c3"),u'(x"10"),u'(x"77"),u'(x"2e"),u'(x"84"),u'(x"83"),
u'(x"82"),u'(x"81"),u'(x"80"),u'(x"87"),u'(x"f7"),u'(x"00"),u'(x"20"),u'(x"0a"),u'(x"f7"),u'(x"00"),u'(x"20"),u'(x"06"),u'(x"f7"),u'(x"00"),u'(x"10"),u'(x"f7"),
u'(x"00"),u'(x"0c"),u'(x"f7"),u'(x"00"),u'(x"04"),u'(x"f7"),u'(x"54"),u'(x"87"),u'(x"26"),u'(x"66"),u'(x"a6"),u'(x"e6"),u'(x"26"),u'(x"66"),u'(x"37"),u'(x"0a"),
u'(x"f7"),u'(x"cc"),u'(x"05"),u'(x"f7"),u'(x"c4"),u'(x"02"),u'(x"77"),u'(x"90"),u'(x"f7"),u'(x"aa"),u'(x"02"),u'(x"10"),u'(x"04"),u'(x"10"),u'(x"f7"),u'(x"24"),
u'(x"7a"),u'(x"f7"),u'(x"76"),u'(x"02"),u'(x"77"),u'(x"74"),u'(x"f7"),u'(x"5e"),u'(x"f7"),u'(x"00"),u'(x"c8"),u'(x"34"),u'(x"f7"),u'(x"6e"),u'(x"74"),u'(x"f7"),
u'(x"7c"),u'(x"70"),u'(x"20"),u'(x"00"),u'(x"00"),u'(x"f7"),u'(x"70"),u'(x"74"),u'(x"10"),u'(x"76"),u'(x"10"),u'(x"f7"),u'(x"5c"),u'(x"4e"),u'(x"f7"),u'(x"5e"),
u'(x"78"),u'(x"10"),u'(x"7a"),u'(x"30"),u'(x"f7"),u'(x"4e"),u'(x"3e"),u'(x"f7"),u'(x"52"),u'(x"c0"),u'(x"34"),u'(x"c0"),u'(x"02"),u'(x"c0"),u'(x"00"),u'(x"02"),
u'(x"c0"),u'(x"fe"),u'(x"37"),u'(x"cc"),u'(x"f7"),u'(x"32"),u'(x"12"),u'(x"20"),u'(x"00"),u'(x"00"),u'(x"f7"),u'(x"26"),u'(x"82"),u'(x"10"),u'(x"00"),u'(x"00"),
u'(x"85"),u'(x"84"),u'(x"83"),u'(x"82"),u'(x"81"),u'(x"80"),u'(x"87"),u'(x"00"),u'(x"22"),u'(x"00"),u'(x"c0"),u'(x"00"),u'(x"c0"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"c0"),u'(x"c0"),u'(x"f7"),u'(x"e0"),u'(x"02"),u'(x"77"),u'(x"80"),u'(x"26"),u'(x"66"),u'(x"a6"),u'(x"e6"),u'(x"26"),u'(x"66"),u'(x"f7"),u'(x"f2"),u'(x"05"),
u'(x"f7"),u'(x"ea"),u'(x"02"),u'(x"77"),u'(x"58"),u'(x"c3"),u'(x"be"),u'(x"37"),u'(x"f4"),u'(x"f7"),u'(x"98"),u'(x"c2"),u'(x"02"),u'(x"c4"),u'(x"00"),u'(x"c4"),
u'(x"fc"),u'(x"c5"),u'(x"f4"),u'(x"37"),u'(x"f6"),u'(x"f7"),u'(x"00"),u'(x"ee"),u'(x"04"),u'(x"f7"),u'(x"00"),u'(x"e6"),u'(x"05"),u'(x"df"),u'(x"00"),u'(x"48"),
u'(x"77"),u'(x"1e"),u'(x"c0"),u'(x"c3"),u'(x"10"),u'(x"02"),u'(x"c0"),u'(x"10"),u'(x"40"),u'(x"01"),u'(x"40"),u'(x"01"),u'(x"c1"),u'(x"01"),u'(x"01"),u'(x"81"),
u'(x"c1"),u'(x"c1"),u'(x"c1"),u'(x"77"),u'(x"0a"),u'(x"f7"),u'(x"70"),u'(x"80"),u'(x"10"),u'(x"60"),u'(x"00"),u'(x"01"),u'(x"c1"),u'(x"01"),u'(x"01"),u'(x"81"),
u'(x"9f"),u'(x"40"),u'(x"1f"),u'(x"42"),u'(x"df"),u'(x"60"),u'(x"44"),u'(x"df"),u'(x"01"),u'(x"47"),u'(x"c1"),u'(x"02"),u'(x"5f"),u'(x"46"),u'(x"01"),u'(x"42"),
u'(x"44"),u'(x"45"),u'(x"77"),u'(x"5e"),u'(x"43"),u'(x"c3"),u'(x"00"),u'(x"38"),u'(x"57"),u'(x"00"),u'(x"33"),u'(x"f7"),u'(x"4e"),u'(x"0a"),u'(x"f7"),u'(x"46"),
u'(x"5e"),u'(x"f7"),u'(x"00"),u'(x"58"),u'(x"f7"),u'(x"00"),u'(x"50"),u'(x"28"),u'(x"f7"),u'(x"00"),u'(x"50"),u'(x"0a"),u'(x"f7"),u'(x"2a"),u'(x"42"),u'(x"f7"),
u'(x"00"),u'(x"3c"),u'(x"f7"),u'(x"00"),u'(x"34"),u'(x"1a"),u'(x"f7"),u'(x"00"),u'(x"2c"),u'(x"f7"),u'(x"34"),u'(x"f7"),u'(x"f8"),u'(x"f2"),u'(x"f7"),u'(x"f4"),
u'(x"ee"),u'(x"f7"),u'(x"a8"),u'(x"c2"),u'(x"12"),u'(x"c4"),u'(x"10"),u'(x"c4"),u'(x"fc"),u'(x"c5"),u'(x"04"),u'(x"37"),u'(x"06"),u'(x"94"),u'(x"77"),u'(x"24"),
u'(x"f7"),u'(x"00"),u'(x"f8"),u'(x"1d"),u'(x"f7"),u'(x"00"),u'(x"f0"),u'(x"f7"),u'(x"00"),u'(x"ea"),u'(x"f7"),u'(x"00"),u'(x"e6"),u'(x"03"),u'(x"f7"),u'(x"c6"),
u'(x"de"),u'(x"f7"),u'(x"c2"),u'(x"03"),u'(x"f7"),u'(x"00"),u'(x"d2"),u'(x"f7"),u'(x"d8"),u'(x"f7"),u'(x"9c"),u'(x"96"),u'(x"f7"),u'(x"98"),u'(x"92"),u'(x"f7"),
u'(x"4c"),u'(x"85"),u'(x"84"),u'(x"83"),u'(x"82"),u'(x"81"),u'(x"80"),u'(x"87"),u'(x"f7"),u'(x"0c"),u'(x"c0"),u'(x"02"),u'(x"77"),u'(x"fe"),u'(x"c0"),u'(x"0a"),
u'(x"f7"),u'(x"5a"),u'(x"02"),u'(x"10"),u'(x"04"),u'(x"10"),u'(x"f7"),u'(x"00"),u'(x"d2"),u'(x"15"),u'(x"f7"),u'(x"64"),u'(x"65"),u'(x"74"),u'(x"74"),u'(x"20"),
u'(x"20"),u'(x"20"),u'(x"20"),u'(x"f7"),u'(x"7a"),u'(x"04"),u'(x"02"),u'(x"f7"),u'(x"4a"),u'(x"0d"),u'(x"00"),u'(x"c0"),u'(x"e3"),u'(x"77"),u'(x"bc"),u'(x"f7"),
u'(x"1c"),u'(x"0a"),u'(x"20"),u'(x"00"),u'(x"00"),u'(x"f7"),u'(x"bc"),u'(x"f7"),u'(x"0c"),u'(x"9a"),u'(x"10"),u'(x"9c"),u'(x"10"),u'(x"f7"),u'(x"1e"),u'(x"1f"),
u'(x"f7"),u'(x"18"),u'(x"69"),u'(x"69"),u'(x"3a"),u'(x"65"),u'(x"64"),u'(x"73"),u'(x"20"),u'(x"69"),u'(x"20"),u'(x"6f"),u'(x"20"),u'(x"65"),u'(x"65"),u'(x"2c"),
u'(x"76"),u'(x"6c"),u'(x"65"),u'(x"69"),u'(x"20"),u'(x"f7"),u'(x"16"),u'(x"9c"),u'(x"02"),u'(x"f7"),u'(x"e6"),u'(x"0d"),u'(x"00"),u'(x"77"),u'(x"5c"),u'(x"f7"),
u'(x"bc"),u'(x"ec"),u'(x"10"),u'(x"fc"),u'(x"30"),u'(x"f7"),u'(x"ce"),u'(x"78"),u'(x"34"),u'(x"36"),u'(x"30"),u'(x"62"),u'(x"61"),u'(x"20"),u'(x"f7"),u'(x"e4"),
u'(x"00"),u'(x"01"),u'(x"f7"),u'(x"b4"),u'(x"3a"),u'(x"f7"),u'(x"d6"),u'(x"01"),u'(x"01"),u'(x"f7"),u'(x"a6"),u'(x"3a"),u'(x"f7"),u'(x"c8"),u'(x"fe"),u'(x"01"),
u'(x"f7"),u'(x"98"),u'(x"3a"),u'(x"f7"),u'(x"ba"),u'(x"ff"),u'(x"01"),u'(x"f7"),u'(x"8a"),u'(x"3a"),u'(x"f7"),u'(x"ac"),u'(x"fc"),u'(x"01"),u'(x"f7"),u'(x"7c"),
u'(x"3a"),u'(x"f7"),u'(x"9e"),u'(x"fd"),u'(x"01"),u'(x"f7"),u'(x"6e"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"ca"),u'(x"40"),u'(x"f7"),u'(x"c5"),u'(x"3b"),u'(x"f7"),
u'(x"bc"),u'(x"36"),u'(x"f7"),u'(x"b7"),u'(x"31"),u'(x"f7"),u'(x"ae"),u'(x"2c"),u'(x"f7"),u'(x"a9"),u'(x"27"),u'(x"f7"),u'(x"00"),u'(x"0e"),u'(x"f7"),u'(x"0a"),
u'(x"ae"),u'(x"f7"),u'(x"18"),u'(x"0e"),u'(x"20"),u'(x"00"),u'(x"00"),u'(x"f7"),u'(x"fe"),u'(x"a0"),u'(x"f7"),u'(x"06"),u'(x"12"),u'(x"20"),u'(x"00"),u'(x"00"),
u'(x"f7"),u'(x"fa"),u'(x"16"),u'(x"10"),u'(x"18"),u'(x"10"),u'(x"f7"),u'(x"0c"),u'(x"65"),u'(x"6f"),u'(x"31"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"f7"),
u'(x"22"),u'(x"18"),u'(x"02"),u'(x"f7"),u'(x"f2"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"cc"),u'(x"1a"),u'(x"20"),u'(x"00"),u'(x"00"),u'(x"f7"),u'(x"c0"),u'(x"16"),
u'(x"10"),u'(x"18"),u'(x"10"),u'(x"f7"),u'(x"d2"),u'(x"65"),u'(x"6f"),u'(x"31"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"f7"),u'(x"e8"),u'(x"18"),u'(x"02"),
u'(x"f7"),u'(x"b8"),u'(x"0d"),u'(x"00"),u'(x"f7"),u'(x"92"),u'(x"22"),u'(x"10"),u'(x"24"),u'(x"10"),u'(x"f7"),u'(x"a4"),u'(x"65"),u'(x"6f"),u'(x"32"),u'(x"20"),
u'(x"20"),u'(x"20"),u'(x"20"),u'(x"f7"),u'(x"ba"),u'(x"24"),u'(x"02"),u'(x"f7"),u'(x"8a"),u'(x"0d"),u'(x"00"),u'(x"00"),u'(x"87"),u'(x"c0"),u'(x"01"),u'(x"87"),
u'(x"c0"),u'(x"0a"),u'(x"f7"),u'(x"52"),u'(x"6e"),u'(x"f7"),u'(x"50"),u'(x"96"),u'(x"20"),u'(x"00"),u'(x"00"),u'(x"37"),u'(x"62"),u'(x"f7"),u'(x"40"),u'(x"9a"),
u'(x"10"),u'(x"9c"),u'(x"10"),u'(x"f7"),u'(x"52"),u'(x"50"),u'(x"22"),u'(x"f7"),u'(x"4a"),u'(x"69"),u'(x"69"),u'(x"3a"),u'(x"65"),u'(x"64"),u'(x"73"),u'(x"20"),
u'(x"69"),u'(x"20"),u'(x"6f"),u'(x"20"),u'(x"65"),u'(x"65"),u'(x"2c"),u'(x"76"),u'(x"6c"),u'(x"65"),u'(x"69"),u'(x"20"),u'(x"f7"),u'(x"48"),u'(x"9c"),u'(x"02"),
u'(x"f7"),u'(x"18"),u'(x"0d"),u'(x"00"),u'(x"c0"),u'(x"cc"),u'(x"c0"),u'(x"01"),u'(x"87"),u'(x"00"),u'(x"87"),u'(x"22"),u'(x"00"),u'(x"20"),u'(x"00"),u'(x"69"),
u'(x"69"),u'(x"3a"),u'(x"65"),u'(x"64"),u'(x"73"),u'(x"20"),u'(x"69"),u'(x"20"),u'(x"6f"),u'(x"20"),u'(x"70"),u'(x"61"),u'(x"65"),u'(x"20"),u'(x"61"),u'(x"75"),
u'(x"20"),u'(x"73"),u'(x"00"),u'(x"6e"),u'(x"74"),u'(x"20"),u'(x"75"),u'(x"61"),u'(x"74"),u'(x"64"),u'(x"64"),u'(x"6e"),u'(x"74"),u'(x"72"),u'(x"73"),u'(x"74"),
u'(x"20"),u'(x"61"),u'(x"75"),u'(x"20"),u'(x"73"),u'(x"00"),u'(x"20"),u'(x"78"),u'(x"34"),u'(x"36"),u'(x"30"),u'(x"62"),u'(x"61"),u'(x"20"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"20"),u'(x"00"),u'(x"20"),u'(x"00"),u'(x"24"),u'(x"10"),u'(x"22"),u'(x"00"),u'(x"22"),u'(x"00"),u'(x"20"),u'(x"00"),u'(x"24"),u'(x"01"),u'(x"24"),
u'(x"02"),u'(x"20"),u'(x"00"),u'(x"24"),u'(x"10"),u'(x"26"),u'(x"10"),u'(x"24"),u'(x"04"),u'(x"26"),u'(x"04"),u'(x"24"),u'(x"02"),u'(x"26"),u'(x"02"),u'(x"f7"),
u'(x"3a"),u'(x"2e"),u'(x"f7"),u'(x"35"),u'(x"29"),u'(x"f7"),u'(x"2c"),u'(x"24"),u'(x"f7"),u'(x"27"),u'(x"1f"),u'(x"f7"),u'(x"1e"),u'(x"1a"),u'(x"f7"),u'(x"19"),
u'(x"15"),u'(x"f7"),u'(x"18"),u'(x"70"),u'(x"40"),u'(x"00"),u'(x"00"),u'(x"87"),u'(x"22"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"66"),
u'(x"85"),u'(x"02"),u'(x"f6"),u'(x"08"),u'(x"02"),u'(x"5f"),u'(x"00"),u'(x"00"),u'(x"5f"),u'(x"04"),u'(x"04"),u'(x"5f"),u'(x"06"),u'(x"06"),u'(x"5f"),u'(x"02"),
u'(x"02"),u'(x"85"),u'(x"87"),u'(x"66"),u'(x"85"),u'(x"02"),u'(x"f6"),u'(x"08"),u'(x"02"),u'(x"5f"),u'(x"00"),u'(x"40"),u'(x"5f"),u'(x"02"),u'(x"42"),u'(x"5f"),
u'(x"04"),u'(x"44"),u'(x"5f"),u'(x"06"),u'(x"46"),u'(x"85"),u'(x"87"),u'(x"df"),u'(x"fc"),u'(x"40"),u'(x"df"),u'(x"f8"),u'(x"42"),u'(x"df"),u'(x"d2"),u'(x"44"),
u'(x"df"),u'(x"00"),u'(x"47"),u'(x"df"),u'(x"08"),u'(x"46"),u'(x"87"),u'(x"df"),u'(x"dc"),u'(x"40"),u'(x"df"),u'(x"d8"),u'(x"42"),u'(x"df"),u'(x"d2"),u'(x"44"),
u'(x"df"),u'(x"01"),u'(x"47"),u'(x"df"),u'(x"08"),u'(x"46"),u'(x"87"),u'(x"df"),u'(x"c2"),u'(x"40"),u'(x"df"),u'(x"be"),u'(x"42"),u'(x"df"),u'(x"1c"),u'(x"44"),
u'(x"df"),u'(x"00"),u'(x"47"),u'(x"df"),u'(x"f0"),u'(x"46"),u'(x"87"),u'(x"df"),u'(x"a2"),u'(x"40"),u'(x"df"),u'(x"9e"),u'(x"42"),u'(x"df"),u'(x"1c"),u'(x"44"),
u'(x"df"),u'(x"01"),u'(x"47"),u'(x"df"),u'(x"d0"),u'(x"46"),u'(x"87"),u'(x"df"),u'(x"3e"),u'(x"40"),u'(x"df"),u'(x"36"),u'(x"42"),u'(x"df"),u'(x"ba"),u'(x"44"),
u'(x"df"),u'(x"00"),u'(x"47"),u'(x"df"),u'(x"08"),u'(x"46"),u'(x"f7"),u'(x"20"),u'(x"18"),u'(x"0b"),u'(x"f7"),u'(x"16"),u'(x"0e"),u'(x"07"),u'(x"f7"),u'(x"00"),
u'(x"10"),u'(x"f7"),u'(x"fc"),u'(x"0c"),u'(x"10"),u'(x"f7"),u'(x"02"),u'(x"04"),u'(x"f7"),u'(x"fa"),u'(x"fc"),u'(x"f7"),u'(x"ea"),u'(x"f8"),u'(x"77"),u'(x"f2"),
u'(x"f7"),u'(x"e0"),u'(x"ee"),u'(x"77"),u'(x"e8"),u'(x"df"),u'(x"e6"),u'(x"40"),u'(x"df"),u'(x"de"),u'(x"42"),u'(x"df"),u'(x"c2"),u'(x"44"),u'(x"df"),u'(x"00"),
u'(x"47"),u'(x"df"),u'(x"08"),u'(x"46"),u'(x"87"),u'(x"26"),u'(x"66"),u'(x"c0"),u'(x"be"),u'(x"c1"),u'(x"b8"),u'(x"c0"),u'(x"04"),u'(x"41"),u'(x"1f"),u'(x"40"),
u'(x"5f"),u'(x"42"),u'(x"df"),u'(x"be"),u'(x"44"),u'(x"df"),u'(x"01"),u'(x"47"),u'(x"df"),u'(x"04"),u'(x"46"),u'(x"f7"),u'(x"01"),u'(x"ce"),u'(x"81"),u'(x"80"),
u'(x"87"),u'(x"26"),u'(x"66"),u'(x"c0"),u'(x"8e"),u'(x"c1"),u'(x"88"),u'(x"c0"),u'(x"04"),u'(x"41"),u'(x"1f"),u'(x"40"),u'(x"5f"),u'(x"42"),u'(x"df"),u'(x"ae"),
u'(x"44"),u'(x"df"),u'(x"01"),u'(x"47"),u'(x"df"),u'(x"04"),u'(x"46"),u'(x"f7"),u'(x"01"),u'(x"98"),u'(x"81"),u'(x"80"),u'(x"87"),u'(x"df"),u'(x"5a"),u'(x"40"),
u'(x"df"),u'(x"52"),u'(x"42"),u'(x"df"),u'(x"aa"),u'(x"44"),u'(x"df"),u'(x"00"),u'(x"47"),u'(x"df"),u'(x"08"),u'(x"46"),u'(x"f7"),u'(x"3c"),u'(x"20"),u'(x"0b"),
u'(x"f7"),u'(x"32"),u'(x"16"),u'(x"07"),u'(x"f7"),u'(x"08"),u'(x"2c"),u'(x"f7"),u'(x"04"),u'(x"28"),u'(x"10"),u'(x"f7"),u'(x"1e"),u'(x"20"),u'(x"f7"),u'(x"16"),
u'(x"18"),u'(x"f7"),u'(x"f2"),u'(x"14"),u'(x"77"),u'(x"0e"),u'(x"f7"),u'(x"e8"),u'(x"0a"),u'(x"77"),u'(x"04"),u'(x"df"),u'(x"02"),u'(x"40"),u'(x"df"),u'(x"fa"),
u'(x"42"),u'(x"df"),u'(x"b2"),u'(x"44"),u'(x"df"),u'(x"00"),u'(x"47"),u'(x"df"),u'(x"08"),u'(x"46"),u'(x"87"),u'(x"26"),u'(x"c0"),u'(x"20"),u'(x"c0"),u'(x"1c"),
u'(x"c0"),u'(x"18"),u'(x"c0"),u'(x"c0"),u'(x"3c"),u'(x"0e"),u'(x"df"),u'(x"04"),u'(x"40"),u'(x"df"),u'(x"00"),u'(x"42"),u'(x"df"),u'(x"de"),u'(x"44"),u'(x"df"),
u'(x"00"),u'(x"47"),u'(x"1f"),u'(x"46"),u'(x"80"),u'(x"87"),u'(x"26"),u'(x"f7"),u'(x"e8"),u'(x"e8"),u'(x"08"),u'(x"c0"),u'(x"e2"),u'(x"c0"),u'(x"de"),u'(x"c0"),
u'(x"da"),u'(x"c0"),u'(x"08"),u'(x"c0"),u'(x"d0"),u'(x"c0"),u'(x"cc"),u'(x"c0"),u'(x"c8"),u'(x"c0"),u'(x"00"),u'(x"c0"),u'(x"3c"),u'(x"0e"),u'(x"df"),u'(x"b4"),
u'(x"40"),u'(x"df"),u'(x"b0"),u'(x"42"),u'(x"df"),u'(x"de"),u'(x"44"),u'(x"df"),u'(x"01"),u'(x"47"),u'(x"1f"),u'(x"46"),u'(x"80"),u'(x"87"),u'(x"f7"),u'(x"04"),
u'(x"30"),u'(x"07"),u'(x"f7"),u'(x"36"),u'(x"26"),u'(x"20"),u'(x"00"),u'(x"00"),u'(x"07"),u'(x"f7"),u'(x"28"),u'(x"2a"),u'(x"20"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"f7"),u'(x"00"),u'(x"0c"),u'(x"07"),u'(x"f7"),u'(x"12"),u'(x"2e"),u'(x"20"),u'(x"00"),u'(x"00"),u'(x"07"),u'(x"f7"),u'(x"04"),u'(x"32"),u'(x"20"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"f7"),u'(x"00"),u'(x"e8"),u'(x"04"),u'(x"f7"),u'(x"01"),u'(x"16"),u'(x"03"),u'(x"37"),u'(x"10"),u'(x"00"),u'(x"87"),u'(x"66"),u'(x"81"),
u'(x"02"),u'(x"df"),u'(x"74"),u'(x"fd"),u'(x"c9"),u'(x"03"),u'(x"5f"),u'(x"76"),u'(x"f8"),u'(x"81"),u'(x"c1"),u'(x"01"),u'(x"01"),u'(x"81"),u'(x"76"),u'(x"02"),
u'(x"81"),u'(x"87"),u'(x"66"),u'(x"85"),u'(x"02"),u'(x"f6"),u'(x"04"),u'(x"02"),u'(x"26"),u'(x"66"),u'(x"a6"),u'(x"42"),u'(x"00"),u'(x"40"),u'(x"02"),u'(x"81"),
u'(x"f7"),u'(x"80"),u'(x"c0"),u'(x"c0"),u'(x"07"),u'(x"df"),u'(x"74"),u'(x"fd"),u'(x"df"),u'(x"20"),u'(x"76"),u'(x"f3"),u'(x"82"),u'(x"81"),u'(x"80"),u'(x"85"),
u'(x"87"),u'(x"66"),u'(x"85"),u'(x"02"),u'(x"f6"),u'(x"04"),u'(x"02"),u'(x"26"),u'(x"66"),u'(x"a6"),u'(x"42"),u'(x"00"),u'(x"40"),u'(x"02"),u'(x"81"),u'(x"c1"),
u'(x"f7"),u'(x"40"),u'(x"c1"),u'(x"f7"),u'(x"3a"),u'(x"c0"),u'(x"c0"),u'(x"0a"),u'(x"c0"),u'(x"c0"),u'(x"07"),u'(x"df"),u'(x"74"),u'(x"fd"),u'(x"df"),u'(x"20"),
u'(x"76"),u'(x"ec"),u'(x"82"),u'(x"81"),u'(x"80"),u'(x"85"),u'(x"87"),u'(x"66"),u'(x"df"),u'(x"74"),u'(x"fd"),u'(x"c9"),u'(x"03"),u'(x"5f"),u'(x"76"),u'(x"f8"),
u'(x"81"),u'(x"87"),u'(x"26"),u'(x"66"),u'(x"40"),u'(x"80"),u'(x"80"),u'(x"80"),u'(x"80"),u'(x"c0"),u'(x"f0"),u'(x"c0"),u'(x"58"),u'(x"df"),u'(x"74"),u'(x"fd"),
u'(x"1f"),u'(x"76"),u'(x"c1"),u'(x"f0"),u'(x"c1"),u'(x"58"),u'(x"df"),u'(x"74"),u'(x"fd"),u'(x"5f"),u'(x"76"),u'(x"81"),u'(x"80"),u'(x"87"),u'(x"26"),u'(x"c0"),
u'(x"02"),u'(x"f7"),u'(x"04"),u'(x"80"),u'(x"87"),u'(x"66"),u'(x"a6"),u'(x"42"),u'(x"81"),u'(x"f7"),u'(x"ae"),u'(x"c0"),u'(x"c0"),u'(x"07"),u'(x"df"),u'(x"74"),
u'(x"fd"),u'(x"df"),u'(x"20"),u'(x"76"),u'(x"f3"),u'(x"82"),u'(x"81"),u'(x"87"),u'(x"37"),u'(x"94"),u'(x"37"),u'(x"94"),u'(x"37"),u'(x"cc"),u'(x"37"),u'(x"92"),
u'(x"37"),u'(x"90"),u'(x"37"),u'(x"8e"),u'(x"37"),u'(x"8c"),u'(x"37"),u'(x"8a"),u'(x"37"),u'(x"8c"),u'(x"37"),u'(x"8a"),u'(x"37"),u'(x"88"),u'(x"37"),u'(x"86"),
u'(x"37"),u'(x"94"),u'(x"37"),u'(x"8e"),u'(x"37"),u'(x"84"),u'(x"37"),u'(x"7e"),u'(x"df"),u'(x"00"),u'(x"48"),u'(x"df"),u'(x"00"),u'(x"4a"),u'(x"df"),u'(x"00"),
u'(x"4c"),u'(x"df"),u'(x"00"),u'(x"4e"),u'(x"87"),u'(x"26"),u'(x"00"),u'(x"80"),u'(x"fe"),u'(x"80"),u'(x"87"),u'(x"b7"),u'(x"36"),u'(x"f7"),u'(x"58"),u'(x"30"),
u'(x"0a"),u'(x"f7"),u'(x"56"),u'(x"64"),u'(x"67"),u'(x"62"),u'(x"72"),u'(x"73"),u'(x"0a"),u'(x"77"),u'(x"aa"),u'(x"02"),u'(x"30"),u'(x"32"),u'(x"34"),u'(x"36"),
u'(x"38"),u'(x"61"),u'(x"63"),u'(x"65"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00") 
);
signal memo : mem_type := mem_type'(
u'(x"00"),u'(x"01"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"15"),u'(x"02"),u'(x"0a"),u'(x"17"),u'(x"15"),u'(x"19"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"09"),u'(x"16"),u'(x"09"),u'(x"17"),u'(x"09"),u'(x"15"),u'(x"65"),u'(x"6c"),u'(x"2c"),u'(x"77"),u'(x"72"),u'(x"64"),u'(x"20"),u'(x"75"),u'(x"63"),u'(x"75"),
u'(x"5b"),u'(x"34"),u'(x"5d"),u'(x"64"),u'(x"75"),u'(x"61"),u'(x"6d"),u'(x"63"),u'(x"6f"),u'(x"6f"),u'(x"65"),u'(x"0a"),u'(x"00"),u'(x"09"),u'(x"0e"),u'(x"0a"),
u'(x"ff"),u'(x"15"),u'(x"08"),u'(x"f9"),u'(x"0b"),u'(x"03"),u'(x"0a"),u'(x"f9"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"f9"),u'(x"01"),u'(x"0a"),u'(x"16"),u'(x"0b"),
u'(x"16"),u'(x"03"),u'(x"09"),u'(x"0c"),u'(x"0b"),u'(x"17"),u'(x"03"),u'(x"55"),u'(x"20"),u'(x"f9"),u'(x"01"),u'(x"0a"),u'(x"11"),u'(x"09"),u'(x"11"),u'(x"14"),
u'(x"00"),u'(x"14"),u'(x"00"),u'(x"0b"),u'(x"11"),u'(x"02"),u'(x"09"),u'(x"14"),u'(x"61"),u'(x"6e"),u'(x"74"),u'(x"72"),u'(x"61"),u'(x"20"),u'(x"69"),u'(x"6c"),
u'(x"64"),u'(x"0a"),u'(x"00"),u'(x"09"),u'(x"0e"),u'(x"09"),u'(x"16"),u'(x"8b"),u'(x"11"),u'(x"02"),u'(x"8b"),u'(x"11"),u'(x"02"),u'(x"8b"),u'(x"11"),u'(x"02"),
u'(x"8b"),u'(x"11"),u'(x"02"),u'(x"8b"),u'(x"11"),u'(x"02"),u'(x"8b"),u'(x"11"),u'(x"03"),u'(x"09"),u'(x"14"),u'(x"65"),u'(x"74"),u'(x"72"),u'(x"6e"),u'(x"20"),
u'(x"61"),u'(x"0d"),u'(x"00"),u'(x"9d"),u'(x"11"),u'(x"11"),u'(x"9d"),u'(x"11"),u'(x"11"),u'(x"9d"),u'(x"11"),u'(x"11"),u'(x"9d"),u'(x"11"),u'(x"11"),u'(x"9d"),
u'(x"11"),u'(x"11"),u'(x"9d"),u'(x"11"),u'(x"11"),u'(x"09"),u'(x"11"),u'(x"0b"),u'(x"16"),u'(x"03"),u'(x"09"),u'(x"14"),u'(x"65"),u'(x"74"),u'(x"72"),u'(x"6e"),
u'(x"20"),u'(x"6f"),u'(x"65"),u'(x"69"),u'(x"73"),u'(x"0a"),u'(x"00"),u'(x"09"),u'(x"13"),u'(x"09"),u'(x"14"),u'(x"68"),u'(x"70"),u'(x"72"),u'(x"73"),u'(x"74"),
u'(x"0a"),u'(x"00"),u'(x"01"),u'(x"09"),u'(x"00"),u'(x"17"),u'(x"f9"),u'(x"45"),u'(x"ff"),u'(x"0b"),u'(x"02"),u'(x"00"),u'(x"ff"),u'(x"25"),u'(x"00"),u'(x"02"),
u'(x"00"),u'(x"fe"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"00"),u'(x"fe"),u'(x"09"),u'(x"14"),u'(x"63"),u'(x"72"),u'(x"20"),u'(x"61"),u'(x"75"),u'(x"20"),u'(x"72"),
u'(x"6e"),u'(x"20"),u'(x"20"),u'(x"00"),u'(x"09"),u'(x"14"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"13"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"fe"),u'(x"17"),u'(x"f9"),
u'(x"35"),u'(x"00"),u'(x"03"),u'(x"8a"),u'(x"f9"),u'(x"00"),u'(x"fe"),u'(x"35"),u'(x"00"),u'(x"02"),u'(x"00"),u'(x"00"),u'(x"8a"),u'(x"f9"),u'(x"45"),u'(x"ff"),
u'(x"10"),u'(x"15"),u'(x"0c"),u'(x"65"),u'(x"05"),u'(x"12"),u'(x"09"),u'(x"00"),u'(x"09"),u'(x"13"),u'(x"63"),u'(x"72"),u'(x"20"),u'(x"6f"),u'(x"70"),u'(x"3a"),
u'(x"00"),u'(x"09"),u'(x"13"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"13"),u'(x"0a"),u'(x"00"),u'(x"55"),u'(x"08"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"13"),u'(x"63"),
u'(x"72"),u'(x"20"),u'(x"6f"),u'(x"70"),u'(x"3a"),u'(x"00"),u'(x"09"),u'(x"13"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"13"),u'(x"0a"),u'(x"00"),u'(x"55"),u'(x"08"),
u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"13"),u'(x"63"),u'(x"72"),u'(x"20"),u'(x"6d"),u'(x"31"),u'(x"67"),u'(x"74"),u'(x"70"),u'(x"62"),u'(x"20"),u'(x"20"),u'(x"00"),
u'(x"09"),u'(x"13"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"13"),u'(x"0a"),u'(x"00"),u'(x"17"),u'(x"f9"),u'(x"15"),u'(x"17"),u'(x"f9"),u'(x"15"),u'(x"55"),u'(x"08"),
u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"13"),u'(x"63"),u'(x"72"),u'(x"20"),u'(x"6d"),u'(x"32"),u'(x"67"),u'(x"74"),u'(x"63"),u'(x"64"),u'(x"20"),u'(x"00"),u'(x"09"),
u'(x"13"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"0a"),u'(x"00"),u'(x"17"),u'(x"f9"),u'(x"00"),u'(x"17"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"0f"),u'(x"00"),
u'(x"00"),u'(x"19"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"63"),u'(x"62"),u'(x"20"),u'(x"6d"),u'(x"32"),u'(x"3a"),u'(x"00"),u'(x"09"),u'(x"13"),u'(x"19"),u'(x"00"),
u'(x"09"),u'(x"12"),u'(x"0a"),u'(x"00"),u'(x"9d"),u'(x"14"),u'(x"a5"),u'(x"00"),u'(x"05"),u'(x"0c"),u'(x"65"),u'(x"05"),u'(x"12"),u'(x"09"),u'(x"00"),u'(x"55"),
u'(x"08"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"63"),u'(x"72"),u'(x"20"),u'(x"54"),u'(x"52"),u'(x"20"),u'(x"20"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"f9"),
u'(x"00"),u'(x"09"),u'(x"12"),u'(x"0a"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"f9"),u'(x"0b"),u'(x"14"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"14"),u'(x"1d"),u'(x"14"),
u'(x"14"),u'(x"1d"),u'(x"14"),u'(x"14"),u'(x"1d"),u'(x"14"),u'(x"14"),u'(x"1d"),u'(x"14"),u'(x"14"),u'(x"55"),u'(x"08"),u'(x"f9"),u'(x"00"),u'(x"55"),u'(x"08"),
u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"07"),u'(x"0b"),u'(x"14"),u'(x"03"),u'(x"55"),u'(x"10"),u'(x"f9"),u'(x"55"),u'(x"08"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"12"),
u'(x"63"),u'(x"72"),u'(x"20"),u'(x"54"),u'(x"50"),u'(x"3a"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"0a"),u'(x"00"),u'(x"0a"),
u'(x"13"),u'(x"15"),u'(x"00"),u'(x"f9"),u'(x"55"),u'(x"08"),u'(x"f9"),u'(x"00"),u'(x"03"),u'(x"04"),u'(x"04"),u'(x"04"),u'(x"05"),u'(x"05"),u'(x"04"),u'(x"04"),
u'(x"05"),u'(x"04"),u'(x"04"),u'(x"04"),u'(x"04"),u'(x"04"),u'(x"04"),u'(x"05"),u'(x"06"),u'(x"06"),u'(x"06"),u'(x"06"),u'(x"07"),u'(x"07"),u'(x"07"),u'(x"08"),
u'(x"09"),u'(x"09"),u'(x"0a"),u'(x"0a"),u'(x"0b"),u'(x"0b"),u'(x"0b"),u'(x"0b"),u'(x"0b"),u'(x"0c"),u'(x"0c"),u'(x"0c"),u'(x"0c"),u'(x"0c"),u'(x"0c"),u'(x"0c"),
u'(x"09"),u'(x"11"),u'(x"63"),u'(x"20"),u'(x"20"),u'(x"6f"),u'(x"70"),u'(x"0a"),u'(x"00"),u'(x"55"),u'(x"08"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"63"),
u'(x"20"),u'(x"20"),u'(x"6f"),u'(x"64"),u'(x"61"),u'(x"64"),u'(x"73"),u'(x"61"),u'(x"74"),u'(x"00"),u'(x"55"),u'(x"40"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"11"),
u'(x"63"),u'(x"20"),u'(x"20"),u'(x"65"),u'(x"64"),u'(x"64"),u'(x"66"),u'(x"75"),u'(x"74"),u'(x"70"),u'(x"79"),u'(x"69"),u'(x"61"),u'(x"20"),u'(x"64"),u'(x"72"),
u'(x"73"),u'(x"20"),u'(x"00"),u'(x"09"),u'(x"0e"),u'(x"09"),u'(x"11"),u'(x"14"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"14"),u'(x"00"),
u'(x"09"),u'(x"11"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"13"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"13"),u'(x"00"),u'(x"09"),u'(x"10"),
u'(x"00"),u'(x"09"),u'(x"11"),u'(x"13"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"13"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"0a"),u'(x"00"),
u'(x"9d"),u'(x"0d"),u'(x"13"),u'(x"9d"),u'(x"0d"),u'(x"13"),u'(x"9d"),u'(x"0d"),u'(x"13"),u'(x"9d"),u'(x"0d"),u'(x"12"),u'(x"9d"),u'(x"0d"),u'(x"12"),u'(x"9d"),
u'(x"0d"),u'(x"12"),u'(x"09"),u'(x"0e"),u'(x"55"),u'(x"08"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"63"),u'(x"20"),u'(x"20"),u'(x"6f"),u'(x"6f"),u'(x"20"),
u'(x"75"),u'(x"63"),u'(x"69"),u'(x"6e"),u'(x"0a"),u'(x"00"),u'(x"55"),u'(x"08"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"63"),u'(x"20"),u'(x"20"),u'(x"65"),
u'(x"64"),u'(x"70"),u'(x"79"),u'(x"69"),u'(x"61"),u'(x"20"),u'(x"64"),u'(x"72"),u'(x"73"),u'(x"20"),u'(x"00"),u'(x"09"),u'(x"0d"),u'(x"9d"),u'(x"0d"),u'(x"12"),
u'(x"9d"),u'(x"0d"),u'(x"12"),u'(x"9d"),u'(x"0d"),u'(x"12"),u'(x"9d"),u'(x"0d"),u'(x"12"),u'(x"9d"),u'(x"0d"),u'(x"12"),u'(x"9d"),u'(x"0d"),u'(x"12"),u'(x"09"),
u'(x"10"),u'(x"19"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"0a"),u'(x"00"),u'(x"09"),u'(x"0d"),u'(x"55"),u'(x"08"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"63"),
u'(x"20"),u'(x"20"),u'(x"72"),u'(x"74"),u'(x"20"),u'(x"68"),u'(x"73"),u'(x"63"),u'(x"6c"),u'(x"61"),u'(x"64"),u'(x"65"),u'(x"73"),u'(x"00"),u'(x"09"),u'(x"0d"),
u'(x"9d"),u'(x"12"),u'(x"0c"),u'(x"9d"),u'(x"12"),u'(x"0c"),u'(x"9d"),u'(x"12"),u'(x"0c"),u'(x"9d"),u'(x"12"),u'(x"0c"),u'(x"9d"),u'(x"12"),u'(x"0c"),u'(x"9d"),
u'(x"12"),u'(x"0c"),u'(x"09"),u'(x"0f"),u'(x"14"),u'(x"00"),u'(x"09"),u'(x"0f"),u'(x"0a"),u'(x"00"),u'(x"09"),u'(x"0c"),u'(x"55"),u'(x"08"),u'(x"f9"),u'(x"00"),
u'(x"09"),u'(x"0f"),u'(x"63"),u'(x"20"),u'(x"20"),u'(x"65"),u'(x"64"),u'(x"6d"),u'(x"6c"),u'(x"69"),u'(x"61"),u'(x"74"),u'(x"61"),u'(x"64"),u'(x"65"),u'(x"73"),
u'(x"6c"),u'(x"73"),u'(x"0d"),u'(x"00"),u'(x"09"),u'(x"0c"),u'(x"9d"),u'(x"11"),u'(x"25"),u'(x"00"),u'(x"05"),u'(x"10"),u'(x"11"),u'(x"0b"),u'(x"03"),u'(x"09"),
u'(x"0e"),u'(x"55"),u'(x"08"),u'(x"f9"),u'(x"00"),u'(x"55"),u'(x"48"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"0f"),u'(x"63"),u'(x"20"),u'(x"20"),u'(x"72"),u'(x"74"),
u'(x"20"),u'(x"75"),u'(x"74"),u'(x"63"),u'(x"73"),u'(x"20"),u'(x"64"),u'(x"72"),u'(x"73"),u'(x"20"),u'(x"69"),u'(x"74"),u'(x"00"),u'(x"09"),u'(x"0c"),u'(x"9d"),
u'(x"11"),u'(x"10"),u'(x"11"),u'(x"0b"),u'(x"02"),u'(x"09"),u'(x"0c"),u'(x"14"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"0f"),u'(x"6c"),u'(x"61"),u'(x"00"),
u'(x"01"),u'(x"25"),u'(x"00"),u'(x"05"),u'(x"09"),u'(x"0b"),u'(x"14"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"0e"),u'(x"09"),u'(x"0f"),u'(x"19"),u'(x"00"),
u'(x"09"),u'(x"0e"),u'(x"0a"),u'(x"00"),u'(x"09"),u'(x"0e"),u'(x"63"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"3a"),u'(x"00"),u'(x"09"),u'(x"0f"),u'(x"19"),
u'(x"00"),u'(x"09"),u'(x"0e"),u'(x"0a"),u'(x"00"),u'(x"09"),u'(x"0e"),u'(x"63"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"3a"),u'(x"00"),u'(x"09"),u'(x"0e"),
u'(x"19"),u'(x"00"),u'(x"09"),u'(x"0e"),u'(x"0a"),u'(x"00"),u'(x"09"),u'(x"0e"),u'(x"63"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"3a"),u'(x"00"),u'(x"09"),
u'(x"0e"),u'(x"19"),u'(x"00"),u'(x"09"),u'(x"0e"),u'(x"0a"),u'(x"00"),u'(x"09"),u'(x"0e"),u'(x"63"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"3a"),u'(x"00"),
u'(x"09"),u'(x"0e"),u'(x"1a"),u'(x"00"),u'(x"09"),u'(x"0e"),u'(x"0a"),u'(x"00"),u'(x"09"),u'(x"0e"),u'(x"63"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"3a"),
u'(x"00"),u'(x"09"),u'(x"0e"),u'(x"1a"),u'(x"00"),u'(x"09"),u'(x"0e"),u'(x"0a"),u'(x"00"),u'(x"55"),u'(x"08"),u'(x"f9"),u'(x"00"),u'(x"55"),u'(x"48"),u'(x"f9"),
u'(x"00"),u'(x"09"),u'(x"0e"),u'(x"63"),u'(x"30"),u'(x"2d"),u'(x"72"),u'(x"61"),u'(x"20"),u'(x"69"),u'(x"67"),u'(x"66"),u'(x"72"),u'(x"61"),u'(x"20"),u'(x"0a"),
u'(x"00"),u'(x"09"),u'(x"0b"),u'(x"1d"),u'(x"0f"),u'(x"10"),u'(x"1d"),u'(x"0f"),u'(x"10"),u'(x"9d"),u'(x"0f"),u'(x"10"),u'(x"1d"),u'(x"0f"),u'(x"10"),u'(x"1d"),
u'(x"0f"),u'(x"10"),u'(x"1d"),u'(x"0f"),u'(x"10"),u'(x"9d"),u'(x"0f"),u'(x"10"),u'(x"1d"),u'(x"0f"),u'(x"10"),u'(x"09"),u'(x"0e"),u'(x"1a"),u'(x"00"),u'(x"09"),
u'(x"0d"),u'(x"0a"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"10"),u'(x"09"),u'(x"0b"),u'(x"55"),u'(x"08"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"0d"),u'(x"63"),u'(x"31"),
u'(x"2d"),u'(x"77"),u'(x"69"),u'(x"65"),u'(x"72"),u'(x"6e"),u'(x"20"),u'(x"6f"),u'(x"6d"),u'(x"74"),u'(x"00"),u'(x"09"),u'(x"0a"),u'(x"15"),u'(x"00"),u'(x"10"),
u'(x"09"),u'(x"0b"),u'(x"09"),u'(x"0d"),u'(x"1a"),u'(x"00"),u'(x"09"),u'(x"0d"),u'(x"0a"),u'(x"00"),u'(x"1d"),u'(x"10"),u'(x"0f"),u'(x"45"),u'(x"00"),u'(x"0f"),
u'(x"1d"),u'(x"0f"),u'(x"0f"),u'(x"45"),u'(x"ff"),u'(x"0f"),u'(x"9d"),u'(x"0f"),u'(x"10"),u'(x"0f"),u'(x"1d"),u'(x"0f"),u'(x"0f"),u'(x"1d"),u'(x"0f"),u'(x"0f"),
u'(x"45"),u'(x"00"),u'(x"0f"),u'(x"1d"),u'(x"0f"),u'(x"0f"),u'(x"45"),u'(x"ff"),u'(x"0f"),u'(x"9d"),u'(x"0f"),u'(x"10"),u'(x"0f"),u'(x"1d"),u'(x"0f"),u'(x"0f"),
u'(x"55"),u'(x"08"),u'(x"f9"),u'(x"1d"),u'(x"0f"),u'(x"0f"),u'(x"1d"),u'(x"0f"),u'(x"0f"),u'(x"1d"),u'(x"0f"),u'(x"0f"),u'(x"1d"),u'(x"0f"),u'(x"0f"),u'(x"1d"),
u'(x"0e"),u'(x"0e"),u'(x"1d"),u'(x"0e"),u'(x"0e"),u'(x"1d"),u'(x"0e"),u'(x"0a"),u'(x"6d"),u'(x"0e"),u'(x"0e"),u'(x"0b"),u'(x"0e"),u'(x"6d"),u'(x"0e"),u'(x"0e"),
u'(x"0b"),u'(x"0e"),u'(x"0a"),u'(x"02"),u'(x"1d"),u'(x"0e"),u'(x"0e"),u'(x"1d"),u'(x"0e"),u'(x"0e"),u'(x"1d"),u'(x"0e"),u'(x"0a"),u'(x"6d"),u'(x"0e"),u'(x"0e"),
u'(x"0b"),u'(x"0e"),u'(x"6d"),u'(x"0e"),u'(x"0e"),u'(x"0b"),u'(x"0e"),u'(x"0a"),u'(x"02"),u'(x"00"),u'(x"09"),u'(x"0c"),u'(x"63"),u'(x"32"),u'(x"2d"),u'(x"72"),
u'(x"61"),u'(x"20"),u'(x"6f"),u'(x"6e"),u'(x"65"),u'(x"73"),u'(x"0a"),u'(x"00"),u'(x"55"),u'(x"08"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"0c"),u'(x"63"),u'(x"33"),
u'(x"2d"),u'(x"72"),u'(x"61"),u'(x"20"),u'(x"6e"),u'(x"20"),u'(x"6c"),u'(x"61"),u'(x"20"),u'(x"6f"),u'(x"6e"),u'(x"65"),u'(x"73"),u'(x"0a"),u'(x"00"),u'(x"55"),
u'(x"08"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"0c"),u'(x"63"),u'(x"34"),u'(x"2d"),u'(x"72"),u'(x"61"),u'(x"20"),u'(x"6f"),u'(x"65"),u'(x"62"),u'(x"74"),u'(x"20"),
u'(x"00"),u'(x"09"),u'(x"0c"),u'(x"19"),u'(x"00"),u'(x"09"),u'(x"0c"),u'(x"0a"),u'(x"00"),u'(x"09"),u'(x"09"),u'(x"1d"),u'(x"0e"),u'(x"0e"),u'(x"09"),u'(x"09"),
u'(x"55"),u'(x"08"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"0c"),u'(x"63"),u'(x"35"),u'(x"2d"),u'(x"77"),u'(x"69"),u'(x"65"),u'(x"6d"),u'(x"64"),u'(x"20"),u'(x"69"),
u'(x"73"),u'(x"00"),u'(x"09"),u'(x"0c"),u'(x"19"),u'(x"00"),u'(x"09"),u'(x"0c"),u'(x"2d"),u'(x"20"),u'(x"00"),u'(x"09"),u'(x"09"),u'(x"1d"),u'(x"0e"),u'(x"0d"),
u'(x"09"),u'(x"0c"),u'(x"19"),u'(x"00"),u'(x"09"),u'(x"0b"),u'(x"0a"),u'(x"00"),u'(x"09"),u'(x"0b"),u'(x"55"),u'(x"08"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"0b"),
u'(x"63"),u'(x"36"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"0b"),u'(x"63"),u'(x"37"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"0b"),u'(x"63"),u'(x"30"),
u'(x"2d"),u'(x"64"),u'(x"6d"),u'(x"20"),u'(x"6e"),u'(x"65"),u'(x"6e"),u'(x"6c"),u'(x"6d"),u'(x"6d"),u'(x"72"),u'(x"0d"),u'(x"00"),u'(x"55"),u'(x"48"),u'(x"f9"),
u'(x"00"),u'(x"09"),u'(x"0b"),u'(x"63"),u'(x"31"),u'(x"2d"),u'(x"6c"),u'(x"61"),u'(x"20"),u'(x"6e"),u'(x"65"),u'(x"6e"),u'(x"6c"),u'(x"6d"),u'(x"6d"),u'(x"72"),
u'(x"0d"),u'(x"00"),u'(x"55"),u'(x"48"),u'(x"f9"),u'(x"00"),u'(x"09"),u'(x"0b"),u'(x"63"),u'(x"32"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"0b"),u'(x"63"),
u'(x"33"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"0b"),u'(x"63"),u'(x"34"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"0b"),u'(x"63"),u'(x"35"),u'(x"0a"),
u'(x"00"),u'(x"00"),u'(x"09"),u'(x"0b"),u'(x"63"),u'(x"36"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"0b"),u'(x"63"),u'(x"37"),u'(x"0a"),u'(x"00"),u'(x"00"),
u'(x"0a"),u'(x"0d"),u'(x"0b"),u'(x"0d"),u'(x"02"),u'(x"0b"),u'(x"0d"),u'(x"02"),u'(x"00"),u'(x"00"),u'(x"10"),u'(x"1d"),u'(x"0c"),u'(x"0d"),u'(x"1d"),u'(x"0c"),
u'(x"0c"),u'(x"0a"),u'(x"0c"),u'(x"09"),u'(x"09"),u'(x"35"),u'(x"80"),u'(x"0c"),u'(x"02"),u'(x"01"),u'(x"0b"),u'(x"0c"),u'(x"03"),u'(x"01"),u'(x"35"),u'(x"02"),
u'(x"0c"),u'(x"02"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"0c"),u'(x"09"),u'(x"00"),u'(x"35"),u'(x"01"),u'(x"0c"),u'(x"03"),u'(x"0a"),u'(x"0c"),u'(x"09"),u'(x"00"),
u'(x"35"),u'(x"01"),u'(x"0c"),u'(x"03"),u'(x"09"),u'(x"00"),u'(x"09"),u'(x"01"),u'(x"2d"),u'(x"0c"),u'(x"0c"),u'(x"02"),u'(x"2d"),u'(x"0c"),u'(x"0c"),u'(x"02"),
u'(x"1d"),u'(x"0c"),u'(x"0c"),u'(x"1d"),u'(x"0c"),u'(x"0c"),u'(x"01"),u'(x"1d"),u'(x"0c"),u'(x"0c"),u'(x"1d"),u'(x"0c"),u'(x"0c"),u'(x"00"),u'(x"ff"),u'(x"15"),
u'(x"00"),u'(x"09"),u'(x"07"),u'(x"0d"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"07"),u'(x"0d"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"0a"),u'(x"0c"),u'(x"00"),
u'(x"88"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"0b"),u'(x"0c"),u'(x"03"),u'(x"55"),u'(x"20"),u'(x"0c"),u'(x"1d"),u'(x"0c"),u'(x"00"),u'(x"09"),u'(x"07"),u'(x"0d"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"07"),u'(x"14"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"07"),u'(x"14"),u'(x"00"),u'(x"14"),u'(x"00"),u'(x"b5"),
u'(x"00"),u'(x"06"),u'(x"02"),u'(x"00"),u'(x"02"),u'(x"00"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"11"),u'(x"1d"),u'(x"0c"),u'(x"1d"),u'(x"0c"),u'(x"45"),
u'(x"00"),u'(x"1d"),u'(x"0c"),u'(x"45"),u'(x"ff"),u'(x"10"),u'(x"25"),u'(x"00"),u'(x"04"),u'(x"15"),u'(x"00"),u'(x"10"),u'(x"35"),u'(x"00"),u'(x"02"),u'(x"01"),
u'(x"0a"),u'(x"10"),u'(x"fe"),u'(x"10"),u'(x"fe"),u'(x"15"),u'(x"1a"),u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"91"),u'(x"fe"),u'(x"0b"),u'(x"0b"),u'(x"02"),
u'(x"0a"),u'(x"0b"),u'(x"ad"),u'(x"06"),u'(x"0c"),u'(x"02"),u'(x"ad"),u'(x"06"),u'(x"0c"),u'(x"02"),u'(x"ad"),u'(x"06"),u'(x"0c"),u'(x"02"),u'(x"ad"),u'(x"06"),
u'(x"0c"),u'(x"02"),u'(x"ad"),u'(x"06"),u'(x"0c"),u'(x"02"),u'(x"ad"),u'(x"06"),u'(x"0c"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"0b"),u'(x"9d"),u'(x"06"),u'(x"0c"),
u'(x"9d"),u'(x"06"),u'(x"0c"),u'(x"9d"),u'(x"06"),u'(x"0c"),u'(x"9d"),u'(x"06"),u'(x"0c"),u'(x"9d"),u'(x"06"),u'(x"0c"),u'(x"9d"),u'(x"06"),u'(x"0c"),u'(x"60"),
u'(x"0b"),u'(x"95"),u'(x"00"),u'(x"0c"),u'(x"95"),u'(x"00"),u'(x"0c"),u'(x"10"),u'(x"0a"),u'(x"0a"),u'(x"0c"),u'(x"0c"),u'(x"0c"),u'(x"11"),u'(x"00"),u'(x"09"),
u'(x"06"),u'(x"1a"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"60"),u'(x"0b"),u'(x"25"),u'(x"00"),u'(x"04"),u'(x"e5"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"15"),u'(x"15"),
u'(x"15"),u'(x"15"),u'(x"15"),u'(x"00"),u'(x"35"),u'(x"01"),u'(x"0b"),u'(x"02"),u'(x"35"),u'(x"80"),u'(x"0b"),u'(x"02"),u'(x"55"),u'(x"40"),u'(x"0b"),u'(x"55"),
u'(x"80"),u'(x"0b"),u'(x"45"),u'(x"80"),u'(x"0b"),u'(x"09"),u'(x"07"),u'(x"00"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"11"),u'(x"11"),u'(x"0a"),u'(x"0b"),
u'(x"0b"),u'(x"0a"),u'(x"02"),u'(x"0b"),u'(x"0a"),u'(x"02"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"05"),u'(x"14"),u'(x"00"),u'(x"14"),u'(x"00"),u'(x"9d"),u'(x"05"),
u'(x"0b"),u'(x"8b"),u'(x"0b"),u'(x"02"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"06"),u'(x"35"),u'(x"80"),u'(x"0a"),u'(x"03"),u'(x"1d"),u'(x"0a"),u'(x"00"),u'(x"09"),
u'(x"05"),u'(x"0f"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"05"),u'(x"0f"),u'(x"00"),u'(x"0f"),u'(x"00"),u'(x"1d"),u'(x"00"),u'(x"0a"),u'(x"09"),u'(x"05"),
u'(x"0f"),u'(x"00"),u'(x"0f"),u'(x"00"),u'(x"1d"),u'(x"00"),u'(x"0a"),u'(x"09"),u'(x"00"),u'(x"1d"),u'(x"0a"),u'(x"e5"),u'(x"00"),u'(x"25"),u'(x"48"),u'(x"05"),
u'(x"15"),u'(x"5f"),u'(x"10"),u'(x"04"),u'(x"09"),u'(x"05"),u'(x"14"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"05"),u'(x"0f"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"15"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"8a"),u'(x"00"),u'(x"2c"),u'(x"00"),u'(x"2c"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"2c"),u'(x"cc"),u'(x"0b"),u'(x"09"),u'(x"02"),u'(x"00"),u'(x"01"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"11"),u'(x"11"),u'(x"0b"),u'(x"09"),u'(x"02"),
u'(x"0b"),u'(x"09"),u'(x"02"),u'(x"00"),u'(x"01"),u'(x"1d"),u'(x"09"),u'(x"0a"),u'(x"09"),u'(x"09"),u'(x"05"),u'(x"1d"),u'(x"0a"),u'(x"1d"),u'(x"0a"),u'(x"45"),
u'(x"ff"),u'(x"1d"),u'(x"09"),u'(x"0a"),u'(x"09"),u'(x"35"),u'(x"80"),u'(x"09"),u'(x"03"),u'(x"55"),u'(x"02"),u'(x"09"),u'(x"01"),u'(x"55"),u'(x"04"),u'(x"f9"),
u'(x"00"),u'(x"01"),u'(x"10"),u'(x"25"),u'(x"00"),u'(x"04"),u'(x"15"),u'(x"00"),u'(x"21"),u'(x"04"),u'(x"11"),u'(x"10"),u'(x"35"),u'(x"00"),u'(x"03"),u'(x"0a"),
u'(x"0c"),u'(x"0c"),u'(x"0c"),u'(x"10"),u'(x"00"),u'(x"09"),u'(x"04"),u'(x"0f"),u'(x"00"),u'(x"1a"),u'(x"00"),u'(x"10"),u'(x"35"),u'(x"00"),u'(x"03"),u'(x"0a"),
u'(x"10"),u'(x"fe"),u'(x"11"),u'(x"fe"),u'(x"15"),u'(x"1a"),u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"0b"),u'(x"03"),u'(x"90"),u'(x"fe"),u'(x"10"),u'(x"60"),
u'(x"0b"),u'(x"e0"),u'(x"60"),u'(x"09"),u'(x"e0"),u'(x"25"),u'(x"00"),u'(x"04"),u'(x"21"),u'(x"00"),u'(x"06"),u'(x"0b"),u'(x"09"),u'(x"03"),u'(x"6d"),u'(x"09"),
u'(x"09"),u'(x"55"),u'(x"80"),u'(x"09"),u'(x"55"),u'(x"40"),u'(x"09"),u'(x"01"),u'(x"35"),u'(x"80"),u'(x"09"),u'(x"02"),u'(x"6d"),u'(x"09"),u'(x"09"),u'(x"55"),
u'(x"80"),u'(x"09"),u'(x"55"),u'(x"40"),u'(x"09"),u'(x"01"),u'(x"45"),u'(x"80"),u'(x"09"),u'(x"09"),u'(x"05"),u'(x"1d"),u'(x"08"),u'(x"08"),u'(x"1d"),u'(x"08"),
u'(x"08"),u'(x"09"),u'(x"04"),u'(x"1d"),u'(x"09"),u'(x"1d"),u'(x"09"),u'(x"45"),u'(x"ff"),u'(x"1d"),u'(x"09"),u'(x"0a"),u'(x"09"),u'(x"01"),u'(x"00"),u'(x"ff"),
u'(x"35"),u'(x"80"),u'(x"08"),u'(x"03"),u'(x"55"),u'(x"01"),u'(x"08"),u'(x"45"),u'(x"80"),u'(x"08"),u'(x"35"),u'(x"80"),u'(x"08"),u'(x"02"),u'(x"6d"),u'(x"08"),
u'(x"08"),u'(x"0b"),u'(x"08"),u'(x"03"),u'(x"55"),u'(x"20"),u'(x"08"),u'(x"09"),u'(x"04"),u'(x"1d"),u'(x"08"),u'(x"08"),u'(x"1d"),u'(x"08"),u'(x"08"),u'(x"09"),
u'(x"04"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"02"),u'(x"0b"),u'(x"03"),u'(x"00"),u'(x"01"),u'(x"15"),u'(x"00"),
u'(x"09"),u'(x"03"),u'(x"14"),u'(x"00"),u'(x"14"),u'(x"00"),u'(x"35"),u'(x"10"),u'(x"02"),u'(x"02"),u'(x"09"),u'(x"06"),u'(x"73"),u'(x"61"),u'(x"20"),u'(x"20"),
u'(x"20"),u'(x"3a"),u'(x"00"),u'(x"09"),u'(x"06"),u'(x"14"),u'(x"00"),u'(x"09"),u'(x"06"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"02"),u'(x"00"),u'(x"01"),u'(x"09"),
u'(x"03"),u'(x"14"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"07"),u'(x"09"),u'(x"03"),u'(x"13"),u'(x"00"),u'(x"13"),u'(x"00"),u'(x"0b"),u'(x"02"),u'(x"03"),
u'(x"09"),u'(x"06"),u'(x"6e"),u'(x"74"),u'(x"20"),u'(x"75"),u'(x"61"),u'(x"74"),u'(x"64"),u'(x"64"),u'(x"6e"),u'(x"74"),u'(x"72"),u'(x"73"),u'(x"74"),u'(x"20"),
u'(x"61"),u'(x"75"),u'(x"20"),u'(x"73"),u'(x"00"),u'(x"09"),u'(x"06"),u'(x"13"),u'(x"00"),u'(x"09"),u'(x"05"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"09"),
u'(x"02"),u'(x"13"),u'(x"00"),u'(x"13"),u'(x"00"),u'(x"09"),u'(x"05"),u'(x"32"),u'(x"6a"),u'(x"30"),u'(x"20"),u'(x"69"),u'(x"3a"),u'(x"00"),u'(x"09"),u'(x"05"),
u'(x"14"),u'(x"00"),u'(x"09"),u'(x"05"),u'(x"00"),u'(x"09"),u'(x"05"),u'(x"14"),u'(x"00"),u'(x"09"),u'(x"05"),u'(x"00"),u'(x"09"),u'(x"05"),u'(x"13"),u'(x"00"),
u'(x"09"),u'(x"05"),u'(x"00"),u'(x"09"),u'(x"05"),u'(x"13"),u'(x"00"),u'(x"09"),u'(x"05"),u'(x"00"),u'(x"09"),u'(x"05"),u'(x"13"),u'(x"00"),u'(x"09"),u'(x"05"),
u'(x"00"),u'(x"09"),u'(x"05"),u'(x"13"),u'(x"00"),u'(x"09"),u'(x"05"),u'(x"0a"),u'(x"00"),u'(x"9d"),u'(x"01"),u'(x"02"),u'(x"9d"),u'(x"01"),u'(x"02"),u'(x"9d"),
u'(x"01"),u'(x"02"),u'(x"9d"),u'(x"01"),u'(x"02"),u'(x"9d"),u'(x"01"),u'(x"02"),u'(x"9d"),u'(x"01"),u'(x"02"),u'(x"15"),u'(x"48"),u'(x"07"),u'(x"1d"),u'(x"07"),
u'(x"01"),u'(x"09"),u'(x"02"),u'(x"14"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"5f"),u'(x"01"),u'(x"09"),u'(x"02"),u'(x"14"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"09"),u'(x"01"),u'(x"14"),u'(x"00"),u'(x"14"),u'(x"00"),u'(x"09"),u'(x"05"),u'(x"63"),u'(x"6e"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"3a"),u'(x"00"),u'(x"09"),
u'(x"05"),u'(x"14"),u'(x"00"),u'(x"09"),u'(x"04"),u'(x"0a"),u'(x"00"),u'(x"09"),u'(x"01"),u'(x"14"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"01"),u'(x"14"),
u'(x"00"),u'(x"14"),u'(x"00"),u'(x"09"),u'(x"04"),u'(x"63"),u'(x"6e"),u'(x"20"),u'(x"20"),u'(x"20"),u'(x"3a"),u'(x"00"),u'(x"09"),u'(x"04"),u'(x"14"),u'(x"00"),
u'(x"09"),u'(x"04"),u'(x"0a"),u'(x"00"),u'(x"09"),u'(x"01"),u'(x"14"),u'(x"00"),u'(x"14"),u'(x"00"),u'(x"09"),u'(x"04"),u'(x"63"),u'(x"6e"),u'(x"20"),u'(x"20"),
u'(x"20"),u'(x"3a"),u'(x"00"),u'(x"09"),u'(x"04"),u'(x"14"),u'(x"00"),u'(x"09"),u'(x"04"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),
u'(x"15"),u'(x"00"),u'(x"15"),u'(x"25"),u'(x"00"),u'(x"09"),u'(x"01"),u'(x"13"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"09"),u'(x"01"),u'(x"13"),
u'(x"00"),u'(x"13"),u'(x"00"),u'(x"25"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"09"),u'(x"04"),u'(x"6e"),u'(x"74"),u'(x"20"),u'(x"75"),u'(x"61"),u'(x"74"),u'(x"64"),
u'(x"64"),u'(x"6e"),u'(x"74"),u'(x"72"),u'(x"73"),u'(x"74"),u'(x"20"),u'(x"61"),u'(x"75"),u'(x"20"),u'(x"73"),u'(x"00"),u'(x"09"),u'(x"04"),u'(x"13"),u'(x"00"),
u'(x"09"),u'(x"04"),u'(x"0a"),u'(x"00"),u'(x"0b"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"36"),u'(x"00"),u'(x"36"),u'(x"00"),u'(x"6e"),
u'(x"74"),u'(x"20"),u'(x"75"),u'(x"61"),u'(x"74"),u'(x"64"),u'(x"64"),u'(x"6e"),u'(x"74"),u'(x"75"),u'(x"64"),u'(x"74"),u'(x"2c"),u'(x"76"),u'(x"6c"),u'(x"65"),
u'(x"69"),u'(x"20"),u'(x"69"),u'(x"69"),u'(x"3a"),u'(x"65"),u'(x"64"),u'(x"73"),u'(x"20"),u'(x"69"),u'(x"20"),u'(x"6f"),u'(x"20"),u'(x"65"),u'(x"65"),u'(x"2c"),
u'(x"76"),u'(x"6c"),u'(x"65"),u'(x"69"),u'(x"20"),u'(x"00"),u'(x"60"),u'(x"32"),u'(x"6a"),u'(x"30"),u'(x"20"),u'(x"69"),u'(x"3a"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"1a"),u'(x"00"),u'(x"74"),u'(x"00"),u'(x"6e"),u'(x"00"),u'(x"04"),u'(x"00"),u'(x"06"),u'(x"00"),u'(x"1e"),u'(x"00"),u'(x"1e"),u'(x"00"),u'(x"1e"),
u'(x"00"),u'(x"6e"),u'(x"00"),u'(x"40"),u'(x"00"),u'(x"40"),u'(x"00"),u'(x"34"),u'(x"00"),u'(x"34"),u'(x"00"),u'(x"34"),u'(x"00"),u'(x"34"),u'(x"00"),u'(x"9d"),
u'(x"00"),u'(x"00"),u'(x"9d"),u'(x"00"),u'(x"00"),u'(x"9d"),u'(x"00"),u'(x"00"),u'(x"9d"),u'(x"00"),u'(x"00"),u'(x"9d"),u'(x"00"),u'(x"00"),u'(x"9d"),u'(x"00"),
u'(x"00"),u'(x"09"),u'(x"00"),u'(x"14"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"60"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"11"),
u'(x"1d"),u'(x"00"),u'(x"65"),u'(x"00"),u'(x"00"),u'(x"1d"),u'(x"00"),u'(x"fe"),u'(x"1d"),u'(x"00"),u'(x"fe"),u'(x"1d"),u'(x"00"),u'(x"fe"),u'(x"1d"),u'(x"00"),
u'(x"fe"),u'(x"15"),u'(x"00"),u'(x"11"),u'(x"1d"),u'(x"00"),u'(x"65"),u'(x"00"),u'(x"00"),u'(x"1d"),u'(x"00"),u'(x"fe"),u'(x"1d"),u'(x"00"),u'(x"fe"),u'(x"1d"),
u'(x"00"),u'(x"fe"),u'(x"1d"),u'(x"00"),u'(x"fe"),u'(x"15"),u'(x"00"),u'(x"1d"),u'(x"04"),u'(x"fe"),u'(x"1d"),u'(x"04"),u'(x"fe"),u'(x"15"),u'(x"19"),u'(x"fe"),
u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"00"),u'(x"1d"),u'(x"04"),u'(x"fe"),u'(x"1d"),u'(x"04"),u'(x"fe"),u'(x"15"),u'(x"19"),u'(x"fe"),
u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"00"),u'(x"1d"),u'(x"04"),u'(x"fe"),u'(x"1d"),u'(x"04"),u'(x"fe"),u'(x"15"),u'(x"1a"),u'(x"fe"),
u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"9d"),u'(x"04"),u'(x"fe"),u'(x"00"),u'(x"1d"),u'(x"04"),u'(x"fe"),u'(x"1d"),u'(x"04"),u'(x"fe"),u'(x"15"),u'(x"1a"),u'(x"fe"),
u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"9d"),u'(x"04"),u'(x"fe"),u'(x"00"),u'(x"1d"),u'(x"04"),u'(x"fe"),u'(x"1d"),u'(x"04"),u'(x"fe"),u'(x"15"),u'(x"19"),u'(x"fe"),
u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"2d"),u'(x"04"),u'(x"04"),u'(x"02"),u'(x"2d"),u'(x"04"),u'(x"04"),u'(x"02"),u'(x"1d"),u'(x"04"),
u'(x"04"),u'(x"1d"),u'(x"03"),u'(x"04"),u'(x"01"),u'(x"1d"),u'(x"04"),u'(x"04"),u'(x"1d"),u'(x"03"),u'(x"03"),u'(x"6d"),u'(x"03"),u'(x"03"),u'(x"0b"),u'(x"03"),
u'(x"6d"),u'(x"03"),u'(x"03"),u'(x"0b"),u'(x"03"),u'(x"1d"),u'(x"03"),u'(x"fe"),u'(x"1d"),u'(x"03"),u'(x"fe"),u'(x"15"),u'(x"19"),u'(x"fe"),u'(x"95"),u'(x"00"),
u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"00"),u'(x"10"),u'(x"10"),u'(x"1d"),u'(x"03"),u'(x"1d"),u'(x"03"),u'(x"65"),u'(x"00"),u'(x"0b"),u'(x"10"),u'(x"fe"),
u'(x"10"),u'(x"fe"),u'(x"15"),u'(x"19"),u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"15"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"15"),
u'(x"00"),u'(x"10"),u'(x"10"),u'(x"1d"),u'(x"03"),u'(x"1d"),u'(x"03"),u'(x"65"),u'(x"00"),u'(x"0b"),u'(x"10"),u'(x"fe"),u'(x"10"),u'(x"fe"),u'(x"15"),u'(x"19"),
u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"15"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"15"),u'(x"00"),u'(x"1d"),u'(x"03"),u'(x"fe"),
u'(x"1d"),u'(x"03"),u'(x"fe"),u'(x"15"),u'(x"19"),u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"2d"),u'(x"03"),u'(x"03"),u'(x"02"),
u'(x"2d"),u'(x"03"),u'(x"03"),u'(x"02"),u'(x"1d"),u'(x"03"),u'(x"03"),u'(x"1d"),u'(x"03"),u'(x"03"),u'(x"01"),u'(x"1d"),u'(x"03"),u'(x"03"),u'(x"1d"),u'(x"03"),
u'(x"03"),u'(x"6d"),u'(x"02"),u'(x"03"),u'(x"0b"),u'(x"03"),u'(x"6d"),u'(x"02"),u'(x"03"),u'(x"0b"),u'(x"03"),u'(x"1d"),u'(x"03"),u'(x"fe"),u'(x"1d"),u'(x"02"),
u'(x"fe"),u'(x"15"),u'(x"19"),u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"00"),u'(x"10"),u'(x"1d"),u'(x"03"),u'(x"6d"),u'(x"03"),
u'(x"6d"),u'(x"03"),u'(x"0c"),u'(x"25"),u'(x"00"),u'(x"05"),u'(x"1d"),u'(x"03"),u'(x"fe"),u'(x"1d"),u'(x"03"),u'(x"fe"),u'(x"15"),u'(x"19"),u'(x"fe"),u'(x"95"),
u'(x"00"),u'(x"fe"),u'(x"90"),u'(x"fe"),u'(x"15"),u'(x"00"),u'(x"10"),u'(x"2d"),u'(x"02"),u'(x"02"),u'(x"06"),u'(x"1d"),u'(x"02"),u'(x"6d"),u'(x"02"),u'(x"6d"),
u'(x"02"),u'(x"0c"),u'(x"01"),u'(x"1d"),u'(x"02"),u'(x"6d"),u'(x"02"),u'(x"6d"),u'(x"02"),u'(x"0c"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"05"),u'(x"1d"),u'(x"02"),
u'(x"fe"),u'(x"1d"),u'(x"02"),u'(x"fe"),u'(x"15"),u'(x"19"),u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"90"),u'(x"fe"),u'(x"15"),u'(x"00"),u'(x"35"),u'(x"00"),
u'(x"02"),u'(x"03"),u'(x"09"),u'(x"fd"),u'(x"14"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"09"),u'(x"fd"),u'(x"14"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"01"),
u'(x"35"),u'(x"80"),u'(x"02"),u'(x"03"),u'(x"09"),u'(x"fd"),u'(x"14"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"09"),u'(x"fd"),u'(x"14"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"01"),u'(x"35"),u'(x"20"),u'(x"01"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"02"),u'(x"01"),u'(x"0a"),u'(x"02"),u'(x"01"),u'(x"00"),u'(x"10"),u'(x"1d"),
u'(x"00"),u'(x"8b"),u'(x"ff"),u'(x"80"),u'(x"8b"),u'(x"03"),u'(x"94"),u'(x"ff"),u'(x"01"),u'(x"0a"),u'(x"35"),u'(x"00"),u'(x"03"),u'(x"0a"),u'(x"10"),u'(x"00"),
u'(x"15"),u'(x"00"),u'(x"11"),u'(x"1d"),u'(x"00"),u'(x"65"),u'(x"00"),u'(x"00"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"1d"),u'(x"00"),u'(x"1d"),u'(x"00"),u'(x"94"),
u'(x"09"),u'(x"00"),u'(x"0a"),u'(x"0b"),u'(x"03"),u'(x"8b"),u'(x"ff"),u'(x"80"),u'(x"95"),u'(x"00"),u'(x"ff"),u'(x"01"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"15"),
u'(x"00"),u'(x"11"),u'(x"1d"),u'(x"00"),u'(x"65"),u'(x"00"),u'(x"00"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"1d"),u'(x"00"),u'(x"1d"),u'(x"00"),u'(x"14"),u'(x"00"),
u'(x"09"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"00"),u'(x"0a"),u'(x"0b"),u'(x"03"),u'(x"0a"),u'(x"0b"),u'(x"03"),u'(x"8b"),u'(x"ff"),u'(x"80"),u'(x"95"),u'(x"00"),
u'(x"ff"),u'(x"01"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"00"),u'(x"10"),u'(x"8b"),u'(x"ff"),u'(x"80"),u'(x"8b"),u'(x"03"),u'(x"94"),u'(x"ff"),u'(x"01"),
u'(x"15"),u'(x"00"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"0c"),u'(x"0c"),u'(x"0c"),u'(x"0c"),u'(x"45"),u'(x"ff"),u'(x"65"),u'(x"19"),u'(x"8b"),u'(x"ff"),u'(x"80"),
u'(x"92"),u'(x"ff"),u'(x"45"),u'(x"ff"),u'(x"65"),u'(x"19"),u'(x"8b"),u'(x"ff"),u'(x"80"),u'(x"92"),u'(x"ff"),u'(x"15"),u'(x"15"),u'(x"00"),u'(x"10"),u'(x"15"),
u'(x"00"),u'(x"09"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"94"),u'(x"09"),u'(x"ff"),u'(x"0a"),u'(x"0b"),u'(x"03"),u'(x"8b"),u'(x"ff"),
u'(x"80"),u'(x"95"),u'(x"00"),u'(x"ff"),u'(x"01"),u'(x"15"),u'(x"15"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"00"),
u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"00"),
u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"f9"),u'(x"15"),u'(x"00"),u'(x"f9"),u'(x"15"),u'(x"00"),
u'(x"f9"),u'(x"15"),u'(x"00"),u'(x"f9"),u'(x"00"),u'(x"10"),u'(x"0a"),u'(x"0a"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"25"),u'(x"02"),u'(x"00"),
u'(x"06"),u'(x"09"),u'(x"fe"),u'(x"6f"),u'(x"20"),u'(x"61"),u'(x"6b"),u'(x"0d"),u'(x"00"),u'(x"00"),u'(x"e8"),u'(x"00"),u'(x"31"),u'(x"33"),u'(x"35"),u'(x"37"),
u'(x"39"),u'(x"62"),u'(x"64"),u'(x"66"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00") 
);


begin
   base_addr_match <= '1' when base_addr(17 downto 13) = bus_addr(17 downto 13) else '0';
   bus_addr_match <= base_addr_match;

   process(clk, base_addr_match)
   begin
      if clk = '1' and clk'event then
         bus_dati(7 downto 0) <= meme(conv_integer(bus_addr(12 downto 1)));
         bus_dati(15 downto 8) <= memo(conv_integer(bus_addr(12 downto 1)));
      end if;
   end process;

   process(clk, base_addr_match)
   begin
      if clk = '1' and clk'event then
         if base_addr_match = '1' and bus_control_dato = '1' then
            if bus_control_datob = '0' or (bus_control_datob = '1' and bus_addr(0) = '0') then
               meme(conv_integer(bus_addr(12 downto 1))) <= bus_dato(7 downto 0);
            end if;
            if bus_control_datob = '0' or (bus_control_datob = '1' and bus_addr(0) = '1') then
               memo(conv_integer(bus_addr(12 downto 1))) <= bus_dato(15 downto 8);
            end if;
         end if;
      end if;
   end process;
end implementation;

