
--
-- Copyright (c) 2008-2020 Sytse van Slooten
--
-- Permission is hereby granted to any person obtaining a copy of these VHDL source files and
-- other language source files and associated documentation files ("the materials") to use
-- these materials solely for personal, non-commercial purposes.
-- You are also granted permission to make changes to the materials, on the condition that this
-- copyright notice is retained unchanged.
--
-- The materials are distributed in the hope that they will be useful, but WITHOUT ANY WARRANTY;
-- without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.
--

-- $Revision$

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity blockram is
   port(
      base_addr : in std_logic_vector(17 downto 0);

      bus_addr_match : out std_logic;
      bus_addr : in std_logic_vector(17 downto 0);
      bus_dati : out std_logic_vector(15 downto 0);
      bus_dato : in std_logic_vector(15 downto 0);
      bus_control_dati : in std_logic;
      bus_control_dato : in std_logic;
      bus_control_datob : in std_logic;

      reset : in std_logic;
      clk : in std_logic
   );
end blockram;

architecture implementation of blockram is

signal base_addr_match : std_logic;

subtype u is std_logic_vector(7 downto 0);
type mem_type is array(0 to 8191) of u;

-- code base at 0

signal meme : mem_type := mem_type'(
u'(x"77"),u'(x"fc"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"c6"),u'(x"fe"),u'(x"77"),u'(x"94"),u'(x"9f"),u'(x"9e"),u'(x"df"),u'(x"9e"),u'(x"78"),u'(x"bf"),u'(x"a4"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"01"),u'(x"78"),
u'(x"00"),u'(x"af"),u'(x"b4"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"02"),u'(x"78"),u'(x"00"),u'(x"af"),u'(x"04"),u'(x"df"),u'(x"03"),u'(x"78"),u'(x"00"),u'(x"b1"),
u'(x"04"),u'(x"df"),u'(x"04"),u'(x"78"),u'(x"00"),u'(x"00"),u'(x"05"),u'(x"08"),u'(x"03"),u'(x"df"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"05"),u'(x"78"),u'(x"00"),
u'(x"df"),u'(x"aa"),u'(x"00"),u'(x"df"),u'(x"aa"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"06"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"55"),u'(x"00"),u'(x"d7"),u'(x"00"),
u'(x"55"),u'(x"04"),u'(x"df"),u'(x"07"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"00"),u'(x"5f"),u'(x"00"),u'(x"d7"),u'(x"00"),u'(x"ff"),u'(x"04"),u'(x"df"),u'(x"08"),
u'(x"78"),u'(x"00"),u'(x"c0"),u'(x"ff"),u'(x"17"),u'(x"ff"),u'(x"04"),u'(x"df"),u'(x"09"),u'(x"78"),u'(x"00"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"04"),u'(x"df"),
u'(x"0a"),u'(x"78"),u'(x"00"),u'(x"c0"),u'(x"aa"),u'(x"17"),u'(x"aa"),u'(x"04"),u'(x"df"),u'(x"0b"),u'(x"78"),u'(x"00"),u'(x"c0"),u'(x"55"),u'(x"17"),u'(x"55"),
u'(x"04"),u'(x"df"),u'(x"0c"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"ff"),u'(x"57"),u'(x"ff"),u'(x"04"),u'(x"df"),u'(x"0d"),u'(x"78"),u'(x"00"),u'(x"01"),u'(x"57"),
u'(x"00"),u'(x"04"),u'(x"df"),u'(x"0e"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"aa"),u'(x"57"),u'(x"aa"),u'(x"04"),u'(x"df"),u'(x"0f"),u'(x"78"),u'(x"00"),u'(x"c1"),
u'(x"55"),u'(x"57"),u'(x"55"),u'(x"04"),u'(x"df"),u'(x"10"),u'(x"78"),u'(x"00"),u'(x"c2"),u'(x"ff"),u'(x"97"),u'(x"ff"),u'(x"04"),u'(x"df"),u'(x"11"),u'(x"78"),
u'(x"00"),u'(x"02"),u'(x"97"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"12"),u'(x"78"),u'(x"00"),u'(x"c2"),u'(x"aa"),u'(x"97"),u'(x"aa"),u'(x"04"),u'(x"df"),u'(x"13"),
u'(x"78"),u'(x"00"),u'(x"c2"),u'(x"55"),u'(x"97"),u'(x"55"),u'(x"04"),u'(x"df"),u'(x"14"),u'(x"78"),u'(x"00"),u'(x"c3"),u'(x"ff"),u'(x"d7"),u'(x"ff"),u'(x"04"),
u'(x"df"),u'(x"15"),u'(x"78"),u'(x"00"),u'(x"03"),u'(x"d7"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"16"),u'(x"78"),u'(x"00"),u'(x"c3"),u'(x"aa"),u'(x"d7"),u'(x"aa"),
u'(x"04"),u'(x"df"),u'(x"17"),u'(x"78"),u'(x"00"),u'(x"c3"),u'(x"55"),u'(x"d7"),u'(x"55"),u'(x"04"),u'(x"df"),u'(x"18"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"ff"),
u'(x"17"),u'(x"ff"),u'(x"04"),u'(x"df"),u'(x"19"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"17"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"1a"),u'(x"78"),u'(x"00"),u'(x"c4"),
u'(x"aa"),u'(x"17"),u'(x"aa"),u'(x"04"),u'(x"df"),u'(x"1b"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"55"),u'(x"17"),u'(x"55"),u'(x"04"),u'(x"df"),u'(x"1c"),u'(x"78"),
u'(x"00"),u'(x"c5"),u'(x"ff"),u'(x"57"),u'(x"ff"),u'(x"04"),u'(x"df"),u'(x"1d"),u'(x"78"),u'(x"00"),u'(x"05"),u'(x"57"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"1e"),
u'(x"78"),u'(x"00"),u'(x"c5"),u'(x"aa"),u'(x"57"),u'(x"aa"),u'(x"04"),u'(x"df"),u'(x"1f"),u'(x"78"),u'(x"00"),u'(x"c5"),u'(x"55"),u'(x"57"),u'(x"55"),u'(x"04"),
u'(x"df"),u'(x"20"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"ff"),u'(x"97"),u'(x"ff"),u'(x"04"),u'(x"df"),u'(x"21"),u'(x"78"),u'(x"00"),u'(x"06"),u'(x"97"),u'(x"00"),
u'(x"04"),u'(x"df"),u'(x"22"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"aa"),u'(x"97"),u'(x"aa"),u'(x"04"),u'(x"df"),u'(x"23"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"55"),
u'(x"97"),u'(x"55"),u'(x"04"),u'(x"df"),u'(x"24"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"ff"),u'(x"fe"),u'(x"df"),u'(x"ef"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"25"),
u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"fe"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"26"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"45"),u'(x"fe"),u'(x"df"),
u'(x"45"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"27"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"aa"),u'(x"fe"),u'(x"df"),u'(x"aa"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"28"),
u'(x"78"),u'(x"00"),u'(x"04"),u'(x"44"),u'(x"04"),u'(x"04"),u'(x"df"),u'(x"29"),u'(x"78"),u'(x"00"),u'(x"44"),u'(x"84"),u'(x"04"),u'(x"df"),u'(x"2a"),u'(x"78"),
u'(x"00"),u'(x"04"),u'(x"44"),u'(x"04"),u'(x"04"),u'(x"df"),u'(x"2b"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"02"),u'(x"44"),u'(x"04"),u'(x"df"),u'(x"2c"),u'(x"78"),
u'(x"00"),u'(x"04"),u'(x"0c"),u'(x"4c"),u'(x"0c"),u'(x"04"),u'(x"df"),u'(x"2d"),u'(x"78"),u'(x"00"),u'(x"4c"),u'(x"03"),u'(x"02"),u'(x"8c"),u'(x"04"),u'(x"df"),
u'(x"2e"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"0c"),u'(x"4c"),u'(x"0c"),u'(x"0c"),u'(x"04"),u'(x"df"),u'(x"2f"),u'(x"78"),u'(x"00"),u'(x"8c"),u'(x"05"),u'(x"04"),
u'(x"4c"),u'(x"8c"),u'(x"8c"),u'(x"04"),u'(x"df"),u'(x"30"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"0c"),u'(x"4c"),u'(x"84"),u'(x"0c"),u'(x"04"),u'(x"df"),u'(x"31"),
u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"8c"),u'(x"84"),u'(x"4c"),u'(x"8c"),u'(x"03"),u'(x"02"),u'(x"8c"),u'(x"04"),u'(x"df"),u'(x"32"),u'(x"78"),u'(x"00"),u'(x"04"),
u'(x"44"),u'(x"84"),u'(x"0c"),u'(x"4c"),u'(x"14"),u'(x"04"),u'(x"df"),u'(x"33"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"c4"),u'(x"54"),u'(x"04"),u'(x"c4"),u'(x"c4"),
u'(x"94"),u'(x"04"),u'(x"df"),u'(x"34"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"44"),u'(x"84"),u'(x"0c"),u'(x"4c"),u'(x"14"),u'(x"04"),u'(x"df"),u'(x"35"),u'(x"78"),
u'(x"00"),u'(x"c4"),u'(x"d4"),u'(x"03"),u'(x"c4"),u'(x"54"),u'(x"04"),u'(x"df"),u'(x"36"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"44"),u'(x"84"),u'(x"0c"),u'(x"4c"),
u'(x"8c"),u'(x"14"),u'(x"04"),u'(x"df"),u'(x"37"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"c4"),u'(x"94"),u'(x"54"),u'(x"03"),u'(x"c4"),u'(x"94"),u'(x"04"),u'(x"df"),
u'(x"38"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"0c"),u'(x"4c"),u'(x"8c"),u'(x"1c"),u'(x"04"),u'(x"df"),u'(x"39"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"c4"),u'(x"5c"),
u'(x"04"),u'(x"c4"),u'(x"c4"),u'(x"9c"),u'(x"04"),u'(x"df"),u'(x"3a"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"01"),u'(x"41"),u'(x"81"),u'(x"09"),u'(x"51"),u'(x"09"),
u'(x"49"),u'(x"0c"),u'(x"4c"),u'(x"8c"),u'(x"1c"),u'(x"04"),u'(x"df"),u'(x"3b"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"c4"),u'(x"5c"),u'(x"c4"),u'(x"c4"),u'(x"9c"),
u'(x"04"),u'(x"df"),u'(x"3c"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"c4"),u'(x"8c"),u'(x"9c"),u'(x"04"),u'(x"c4"),u'(x"c4"),u'(x"1c"),u'(x"04"),u'(x"df"),u'(x"3d"),
u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"c4"),u'(x"5c"),u'(x"c4"),u'(x"c4"),u'(x"9c"),u'(x"04"),u'(x"df"),u'(x"3e"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"44"),u'(x"84"),
u'(x"0c"),u'(x"54"),u'(x"0c"),u'(x"94"),u'(x"24"),u'(x"04"),u'(x"df"),u'(x"3f"),u'(x"78"),u'(x"00"),u'(x"e4"),u'(x"4c"),u'(x"05"),u'(x"04"),u'(x"84"),u'(x"84"),
u'(x"e4"),u'(x"04"),u'(x"df"),u'(x"40"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"44"),u'(x"84"),u'(x"24"),u'(x"4c"),u'(x"94"),u'(x"0c"),u'(x"54"),u'(x"84"),u'(x"24"),
u'(x"04"),u'(x"df"),u'(x"41"),u'(x"78"),u'(x"00"),u'(x"84"),u'(x"84"),u'(x"64"),u'(x"c4"),u'(x"c4"),u'(x"a4"),u'(x"04"),u'(x"df"),u'(x"42"),u'(x"78"),u'(x"00"),
u'(x"e4"),u'(x"04"),u'(x"df"),u'(x"43"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"0c"),u'(x"4c"),u'(x"94"),u'(x"2c"),u'(x"04"),u'(x"df"),u'(x"44"),u'(x"78"),u'(x"00"),
u'(x"84"),u'(x"84"),u'(x"6c"),u'(x"07"),u'(x"84"),u'(x"84"),u'(x"ec"),u'(x"03"),u'(x"94"),u'(x"ac"),u'(x"04"),u'(x"df"),u'(x"45"),u'(x"78"),u'(x"00"),u'(x"04"),
u'(x"44"),u'(x"84"),u'(x"01"),u'(x"41"),u'(x"c1"),u'(x"02"),u'(x"0a"),u'(x"0c"),u'(x"4c"),u'(x"09"),u'(x"2c"),u'(x"04"),u'(x"df"),u'(x"46"),u'(x"78"),u'(x"00"),
u'(x"dc"),u'(x"2c"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"47"),u'(x"78"),u'(x"00"),u'(x"dc"),u'(x"04"),u'(x"df"),u'(x"48"),u'(x"78"),u'(x"00"),
u'(x"8a"),u'(x"2c"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"49"),u'(x"78"),u'(x"00"),u'(x"8a"),u'(x"04"),u'(x"df"),u'(x"4a"),u'(x"78"),u'(x"00"),
u'(x"04"),u'(x"84"),u'(x"84"),u'(x"01"),u'(x"41"),u'(x"81"),u'(x"09"),u'(x"51"),u'(x"09"),u'(x"89"),u'(x"02"),u'(x"0a"),u'(x"34"),u'(x"fe"),u'(x"04"),u'(x"df"),
u'(x"4b"),u'(x"78"),u'(x"00"),u'(x"f4"),u'(x"fe"),u'(x"74"),u'(x"00"),u'(x"05"),u'(x"b4"),u'(x"00"),u'(x"b4"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"4c"),u'(x"78"),
u'(x"00"),u'(x"b1"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"4d"),u'(x"78"),u'(x"00"),u'(x"01"),u'(x"04"),u'(x"44"),u'(x"84"),u'(x"0c"),u'(x"4c"),u'(x"24"),u'(x"24"),
u'(x"94"),u'(x"34"),u'(x"02"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"4e"),u'(x"78"),u'(x"00"),u'(x"f4"),u'(x"02"),u'(x"04"),u'(x"df"),u'(x"4f"),
u'(x"78"),u'(x"00"),u'(x"34"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"50"),u'(x"78"),u'(x"00"),u'(x"31"),u'(x"fc"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),
u'(x"51"),u'(x"78"),u'(x"00"),u'(x"b1"),u'(x"fc"),u'(x"04"),u'(x"df"),u'(x"52"),u'(x"78"),u'(x"00"),u'(x"01"),u'(x"04"),u'(x"44"),u'(x"84"),u'(x"09"),u'(x"49"),
u'(x"89"),u'(x"89"),u'(x"89"),u'(x"0c"),u'(x"34"),u'(x"02"),u'(x"74"),u'(x"02"),u'(x"3c"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"53"),u'(x"78"),u'(x"00"),u'(x"79"),
u'(x"00"),u'(x"04"),u'(x"df"),u'(x"54"),u'(x"78"),u'(x"00"),u'(x"44"),u'(x"bc"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"55"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"0c"),
u'(x"02"),u'(x"42"),u'(x"82"),u'(x"0a"),u'(x"3a"),u'(x"00"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"56"),u'(x"78"),u'(x"00"),u'(x"cc"),u'(x"3c"),u'(x"00"),u'(x"03"),
u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"57"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"44"),u'(x"84"),u'(x"17"),u'(x"ff"),u'(x"04"),u'(x"df"),u'(x"58"),u'(x"78"),
u'(x"00"),u'(x"04"),u'(x"bf"),u'(x"a4"),u'(x"c4"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"59"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"bf"),u'(x"a8"),
u'(x"c4"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"5a"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"44"),u'(x"bf"),u'(x"a8"),u'(x"c4"),u'(x"03"),u'(x"02"),
u'(x"01"),u'(x"04"),u'(x"df"),u'(x"5b"),u'(x"78"),u'(x"00"),u'(x"84"),u'(x"c4"),u'(x"04"),u'(x"df"),u'(x"5c"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"0c"),u'(x"bf"),
u'(x"a4"),u'(x"cc"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"5d"),u'(x"78"),u'(x"00"),u'(x"8c"),u'(x"bf"),u'(x"cc"),u'(x"03"),u'(x"02"),u'(x"01"),
u'(x"04"),u'(x"df"),u'(x"5e"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"0c"),u'(x"4c"),u'(x"8c"),u'(x"bf"),u'(x"a4"),u'(x"cc"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),
u'(x"df"),u'(x"5f"),u'(x"78"),u'(x"00"),u'(x"84"),u'(x"bf"),u'(x"cc"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"60"),u'(x"78"),u'(x"00"),u'(x"04"),
u'(x"14"),u'(x"0c"),u'(x"4c"),u'(x"04"),u'(x"bf"),u'(x"a4"),u'(x"d4"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"61"),u'(x"78"),u'(x"00"),u'(x"d4"),
u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"62"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"14"),u'(x"64"),u'(x"c4"),u'(x"bf"),u'(x"a4"),u'(x"d4"),u'(x"03"),
u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"63"),u'(x"78"),u'(x"00"),u'(x"bf"),u'(x"a8"),u'(x"d4"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"64"),
u'(x"78"),u'(x"00"),u'(x"04"),u'(x"0c"),u'(x"4c"),u'(x"8c"),u'(x"1c"),u'(x"04"),u'(x"bf"),u'(x"a4"),u'(x"dc"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),
u'(x"65"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"c4"),u'(x"dc"),u'(x"04"),u'(x"bf"),u'(x"a8"),u'(x"dc"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"66"),
u'(x"78"),u'(x"00"),u'(x"04"),u'(x"0c"),u'(x"4c"),u'(x"8c"),u'(x"01"),u'(x"41"),u'(x"81"),u'(x"09"),u'(x"bf"),u'(x"dc"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),
u'(x"df"),u'(x"67"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"c4"),u'(x"c4"),u'(x"04"),u'(x"df"),u'(x"68"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"0c"),u'(x"4c"),u'(x"8c"),
u'(x"8c"),u'(x"01"),u'(x"41"),u'(x"81"),u'(x"09"),u'(x"49"),u'(x"09"),u'(x"dc"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"69"),u'(x"78"),u'(x"00"),
u'(x"c4"),u'(x"c4"),u'(x"04"),u'(x"df"),u'(x"6a"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"0c"),u'(x"84"),u'(x"84"),u'(x"bf"),u'(x"a4"),u'(x"e4"),u'(x"03"),u'(x"02"),
u'(x"01"),u'(x"04"),u'(x"df"),u'(x"6b"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"04"),u'(x"df"),u'(x"6c"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"0c"),u'(x"4c"),u'(x"4c"),
u'(x"bf"),u'(x"84"),u'(x"84"),u'(x"e4"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"6d"),u'(x"78"),u'(x"00"),u'(x"e4"),u'(x"04"),u'(x"df"),u'(x"6e"),
u'(x"78"),u'(x"00"),u'(x"04"),u'(x"14"),u'(x"bf"),u'(x"a4"),u'(x"ec"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"6f"),u'(x"78"),u'(x"00"),u'(x"c4"),
u'(x"04"),u'(x"df"),u'(x"70"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"0c"),u'(x"4c"),u'(x"8c"),u'(x"1c"),u'(x"6c"),u'(x"5c"),u'(x"ec"),u'(x"03"),u'(x"02"),u'(x"01"),
u'(x"04"),u'(x"df"),u'(x"71"),u'(x"78"),u'(x"00"),u'(x"94"),u'(x"ec"),u'(x"04"),u'(x"df"),u'(x"72"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"0c"),u'(x"44"),u'(x"84"),
u'(x"0c"),u'(x"4c"),u'(x"f4"),u'(x"00"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"73"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"f4"),u'(x"00"),u'(x"01"),
u'(x"04"),u'(x"df"),u'(x"74"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"0c"),u'(x"54"),u'(x"0c"),u'(x"02"),u'(x"04"),u'(x"44"),u'(x"84"),u'(x"0c"),u'(x"fc"),u'(x"02"),
u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"75"),u'(x"78"),u'(x"00"),u'(x"92"),u'(x"fc"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"76"),u'(x"78"),
u'(x"00"),u'(x"04"),u'(x"01"),u'(x"41"),u'(x"44"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"77"),u'(x"78"),u'(x"00"),u'(x"84"),u'(x"fa"),u'(x"04"),u'(x"01"),
u'(x"41"),u'(x"44"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"78"),u'(x"78"),u'(x"00"),u'(x"84"),u'(x"04"),u'(x"df"),u'(x"79"),u'(x"78"),u'(x"00"),
u'(x"04"),u'(x"01"),u'(x"81"),u'(x"44"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"7a"),u'(x"78"),u'(x"00"),u'(x"41"),u'(x"81"),u'(x"44"),u'(x"04"),
u'(x"df"),u'(x"7b"),u'(x"78"),u'(x"00"),u'(x"af"),u'(x"c4"),u'(x"aa"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"7c"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"55"),u'(x"01"),
u'(x"04"),u'(x"df"),u'(x"7d"),u'(x"78"),u'(x"00"),u'(x"44"),u'(x"04"),u'(x"df"),u'(x"7e"),u'(x"78"),u'(x"00"),u'(x"84"),u'(x"fa"),u'(x"04"),u'(x"44"),u'(x"c1"),
u'(x"aa"),u'(x"c2"),u'(x"55"),u'(x"b1"),u'(x"44"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"7f"),u'(x"78"),u'(x"00"),u'(x"02"),u'(x"04"),u'(x"df"),
u'(x"80"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"81"),u'(x"04"),u'(x"df"),u'(x"81"),u'(x"78"),u'(x"00"),u'(x"81"),u'(x"81"),u'(x"81"),u'(x"f8"),u'(x"c1"),u'(x"aa"),
u'(x"c4"),u'(x"00"),u'(x"c2"),u'(x"55"),u'(x"01"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"82"),u'(x"78"),u'(x"00"),u'(x"01"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),
u'(x"83"),u'(x"78"),u'(x"00"),u'(x"44"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"84"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"84"),u'(x"bf"),u'(x"01"),
u'(x"04"),u'(x"df"),u'(x"85"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"00"),u'(x"c1"),u'(x"02"),u'(x"0c"),u'(x"4c"),u'(x"09"),u'(x"49"),u'(x"02"),u'(x"c3"),u'(x"05"),
u'(x"bf"),u'(x"0a"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"86"),u'(x"78"),u'(x"00"),u'(x"8a"),u'(x"04"),u'(x"af"),u'(x"4b"),u'(x"01"),u'(x"04"),
u'(x"df"),u'(x"87"),u'(x"78"),u'(x"00"),u'(x"8b"),u'(x"fa"),u'(x"02"),u'(x"42"),u'(x"05"),u'(x"04"),u'(x"03"),u'(x"c2"),u'(x"ff"),u'(x"04"),u'(x"df"),u'(x"88"),
u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"00"),u'(x"c1"),u'(x"02"),u'(x"cc"),u'(x"eb"),u'(x"c9"),u'(x"14"),u'(x"4c"),u'(x"04"),u'(x"03"),u'(x"02"),u'(x"8c"),u'(x"04"),
u'(x"df"),u'(x"89"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"00"),u'(x"c1"),u'(x"04"),u'(x"cc"),u'(x"03"),u'(x"c9"),u'(x"06"),u'(x"bf"),u'(x"09"),u'(x"02"),u'(x"01"),
u'(x"04"),u'(x"df"),u'(x"8a"),u'(x"78"),u'(x"00"),u'(x"09"),u'(x"fa"),u'(x"c4"),u'(x"00"),u'(x"c1"),u'(x"02"),u'(x"cc"),u'(x"55"),u'(x"c9"),u'(x"aa"),u'(x"09"),
u'(x"01"),u'(x"04"),u'(x"df"),u'(x"8b"),u'(x"78"),u'(x"00"),u'(x"89"),u'(x"04"),u'(x"df"),u'(x"8c"),u'(x"78"),u'(x"00"),u'(x"c9"),u'(x"09"),u'(x"01"),u'(x"04"),
u'(x"df"),u'(x"8d"),u'(x"78"),u'(x"00"),u'(x"49"),u'(x"4c"),u'(x"04"),u'(x"df"),u'(x"8e"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"00"),u'(x"cc"),u'(x"55"),u'(x"c1"),
u'(x"02"),u'(x"c9"),u'(x"aa"),u'(x"a1"),u'(x"09"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"8f"),u'(x"78"),u'(x"00"),u'(x"09"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),
u'(x"df"),u'(x"90"),u'(x"78"),u'(x"00"),u'(x"0c"),u'(x"8c"),u'(x"4c"),u'(x"04"),u'(x"df"),u'(x"91"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"00"),u'(x"c1"),u'(x"02"),
u'(x"cc"),u'(x"05"),u'(x"11"),u'(x"09"),u'(x"49"),u'(x"e1"),u'(x"bf"),u'(x"54"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"92"),u'(x"78"),u'(x"00"),
u'(x"a4"),u'(x"09"),u'(x"04"),u'(x"df"),u'(x"93"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"00"),u'(x"c1"),u'(x"02"),u'(x"cc"),u'(x"f0"),u'(x"c9"),u'(x"e8"),u'(x"11"),
u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"94"),u'(x"78"),u'(x"00"),u'(x"a1"),u'(x"d1"),u'(x"f9"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"95"),u'(x"78"),
u'(x"00"),u'(x"c4"),u'(x"00"),u'(x"c1"),u'(x"02"),u'(x"c2"),u'(x"04"),u'(x"cc"),u'(x"01"),u'(x"c9"),u'(x"05"),u'(x"d2"),u'(x"38"),u'(x"d2"),u'(x"ff"),u'(x"11"),
u'(x"01"),u'(x"04"),u'(x"df"),u'(x"96"),u'(x"78"),u'(x"00"),u'(x"11"),u'(x"11"),u'(x"c1"),u'(x"11"),u'(x"04"),u'(x"df"),u'(x"97"),u'(x"78"),u'(x"00"),u'(x"8c"),
u'(x"04"),u'(x"df"),u'(x"98"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"00"),u'(x"c1"),u'(x"02"),u'(x"cc"),u'(x"aa"),u'(x"d1"),u'(x"01"),u'(x"c9"),u'(x"02"),u'(x"e1"),
u'(x"11"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"99"),u'(x"78"),u'(x"00"),u'(x"54"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"9a"),u'(x"78"),u'(x"00"),u'(x"11"),u'(x"02"),
u'(x"01"),u'(x"04"),u'(x"df"),u'(x"9b"),u'(x"78"),u'(x"00"),u'(x"e1"),u'(x"e1"),u'(x"54"),u'(x"04"),u'(x"df"),u'(x"9c"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"c1"),
u'(x"02"),u'(x"c2"),u'(x"00"),u'(x"cc"),u'(x"00"),u'(x"c9"),u'(x"02"),u'(x"d2"),u'(x"80"),u'(x"ca"),u'(x"d0"),u'(x"19"),u'(x"00"),u'(x"02"),u'(x"01"),u'(x"04"),
u'(x"df"),u'(x"9d"),u'(x"78"),u'(x"00"),u'(x"ca"),u'(x"50"),u'(x"04"),u'(x"df"),u'(x"9e"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"00"),u'(x"c1"),u'(x"02"),u'(x"d1"),
u'(x"f6"),u'(x"d4"),u'(x"01"),u'(x"21"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"9f"),u'(x"78"),u'(x"00"),u'(x"84"),u'(x"81"),u'(x"b1"),u'(x"64"),u'(x"01"),u'(x"04"),
u'(x"df"),u'(x"a0"),u'(x"78"),u'(x"00"),u'(x"d4"),u'(x"81"),u'(x"21"),u'(x"04"),u'(x"df"),u'(x"a1"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"00"),u'(x"d4"),u'(x"01"),
u'(x"d4"),u'(x"fe"),u'(x"d4"),u'(x"00"),u'(x"cc"),u'(x"02"),u'(x"c1"),u'(x"08"),u'(x"29"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"a2"),u'(x"78"),u'(x"00"),
u'(x"c4"),u'(x"04"),u'(x"6c"),u'(x"04"),u'(x"df"),u'(x"a3"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"c1"),u'(x"00"),u'(x"d1"),u'(x"aa"),u'(x"d1"),u'(x"01"),u'(x"d1"),
u'(x"00"),u'(x"31"),u'(x"00"),u'(x"fc"),u'(x"04"),u'(x"df"),u'(x"a4"),u'(x"78"),u'(x"00"),u'(x"31"),u'(x"05"),u'(x"fa"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"a5"),
u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"00"),u'(x"01"),u'(x"d4"),u'(x"fe"),u'(x"d4"),u'(x"ff"),u'(x"d4"),u'(x"00"),u'(x"c9"),u'(x"02"),u'(x"81"),u'(x"39"),u'(x"fa"),
u'(x"03"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"a6"),u'(x"78"),u'(x"00"),u'(x"7c"),u'(x"ff"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"a7"),u'(x"78"),u'(x"00"),u'(x"c4"),
u'(x"aa"),u'(x"bf"),u'(x"44"),u'(x"04"),u'(x"03"),u'(x"c4"),u'(x"55"),u'(x"04"),u'(x"df"),u'(x"a8"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"aa"),u'(x"af"),u'(x"44"),
u'(x"05"),u'(x"04"),u'(x"03"),u'(x"c4"),u'(x"54"),u'(x"04"),u'(x"df"),u'(x"a9"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"cc"),u'(x"55"),u'(x"4c"),u'(x"05"),u'(x"04"),
u'(x"03"),u'(x"17"),u'(x"aa"),u'(x"04"),u'(x"df"),u'(x"aa"),u'(x"78"),u'(x"00"),u'(x"cc"),u'(x"aa"),u'(x"84"),u'(x"bf"),u'(x"4c"),u'(x"06"),u'(x"05"),u'(x"04"),
u'(x"c4"),u'(x"cc"),u'(x"aa"),u'(x"04"),u'(x"df"),u'(x"ab"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"cc"),u'(x"00"),u'(x"af"),u'(x"54"),u'(x"02"),u'(x"01"),u'(x"04"),
u'(x"df"),u'(x"ac"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"c4"),u'(x"0a"),u'(x"cc"),u'(x"20"),u'(x"a1"),u'(x"54"),u'(x"05"),u'(x"04"),u'(x"c4"),u'(x"cc"),u'(x"40"),
u'(x"04"),u'(x"df"),u'(x"ad"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"cc"),u'(x"55"),u'(x"bf"),u'(x"5f"),u'(x"00"),u'(x"05"),u'(x"04"),u'(x"03"),u'(x"cc"),u'(x"ab"),
u'(x"04"),u'(x"df"),u'(x"ae"),u'(x"78"),u'(x"00"),u'(x"cc"),u'(x"aa"),u'(x"b1"),u'(x"5f"),u'(x"00"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"af"),u'(x"78"),
u'(x"00"),u'(x"01"),u'(x"c4"),u'(x"02"),u'(x"c9"),u'(x"d1"),u'(x"bf"),u'(x"64"),u'(x"07"),u'(x"06"),u'(x"05"),u'(x"c9"),u'(x"a3"),u'(x"02"),u'(x"c4"),u'(x"04"),
u'(x"df"),u'(x"b0"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"cc"),u'(x"00"),u'(x"dc"),u'(x"2e"),u'(x"bf"),u'(x"6c"),u'(x"08"),u'(x"07"),u'(x"06"),u'(x"c4"),u'(x"04"),
u'(x"df"),u'(x"5d"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"b1"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"00"),u'(x"01"),u'(x"c9"),u'(x"55"),u'(x"bf"),u'(x"74"),u'(x"00"),
u'(x"05"),u'(x"04"),u'(x"03"),u'(x"c9"),u'(x"ab"),u'(x"04"),u'(x"df"),u'(x"b2"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"00"),u'(x"1f"),u'(x"02"),u'(x"df"),u'(x"00"),
u'(x"00"),u'(x"7c"),u'(x"02"),u'(x"06"),u'(x"05"),u'(x"04"),u'(x"03"),u'(x"df"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"b3"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"00"),
u'(x"cc"),u'(x"c0"),u'(x"df"),u'(x"00"),u'(x"06"),u'(x"cc"),u'(x"41"),u'(x"03"),u'(x"df"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"b4"),u'(x"78"),u'(x"00"),u'(x"c4"),
u'(x"55"),u'(x"af"),u'(x"04"),u'(x"03"),u'(x"c4"),u'(x"aa"),u'(x"04"),u'(x"df"),u'(x"b5"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"cc"),u'(x"01"),u'(x"bf"),u'(x"0c"),
u'(x"04"),u'(x"03"),u'(x"cc"),u'(x"80"),u'(x"04"),u'(x"df"),u'(x"b6"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"01"),u'(x"cc"),u'(x"c1"),u'(x"68"),u'(x"49"),u'(x"d7"),
u'(x"cc"),u'(x"02"),u'(x"04"),u'(x"df"),u'(x"b7"),u'(x"78"),u'(x"00"),u'(x"57"),u'(x"40"),u'(x"04"),u'(x"df"),u'(x"b8"),u'(x"78"),u'(x"00"),u'(x"9f"),u'(x"cc"),
u'(x"c1"),u'(x"66"),u'(x"59"),u'(x"82"),u'(x"d7"),u'(x"cc"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"b9"),u'(x"78"),u'(x"00"),u'(x"9f"),u'(x"cc"),u'(x"c1"),u'(x"3e"),
u'(x"51"),u'(x"d7"),u'(x"cc"),u'(x"03"),u'(x"04"),u'(x"df"),u'(x"ba"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"68"),u'(x"04"),u'(x"df"),u'(x"bb"),u'(x"78"),u'(x"00"),
u'(x"9f"),u'(x"cc"),u'(x"c1"),u'(x"d8"),u'(x"61"),u'(x"00"),u'(x"c1"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"bc"),u'(x"78"),u'(x"00"),u'(x"d7"),u'(x"cc"),u'(x"05"),
u'(x"04"),u'(x"df"),u'(x"bd"),u'(x"78"),u'(x"00"),u'(x"9f"),u'(x"cc"),u'(x"c1"),u'(x"fd"),u'(x"71"),u'(x"05"),u'(x"a0"),u'(x"c1"),u'(x"d6"),u'(x"04"),u'(x"df"),
u'(x"be"),u'(x"78"),u'(x"00"),u'(x"d7"),u'(x"cc"),u'(x"04"),u'(x"04"),u'(x"df"),u'(x"bf"),u'(x"78"),u'(x"00"),u'(x"9f"),u'(x"cc"),u'(x"c1"),u'(x"02"),u'(x"69"),
u'(x"ac"),u'(x"df"),u'(x"06"),u'(x"cc"),u'(x"04"),u'(x"df"),u'(x"c0"),u'(x"78"),u'(x"00"),u'(x"9f"),u'(x"cc"),u'(x"c1"),u'(x"26"),u'(x"79"),u'(x"f8"),u'(x"22"),
u'(x"00"),u'(x"df"),u'(x"07"),u'(x"cc"),u'(x"04"),u'(x"df"),u'(x"c1"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"fa"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),
u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),
u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),
u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),
u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),
u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),
u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"cf"),u'(x"a0"),u'(x"49"),u'(x"5f"),u'(x"02"),u'(x"df"),u'(x"c2"),u'(x"78"),
u'(x"00"),u'(x"c2"),u'(x"20"),u'(x"c3"),u'(x"3a"),u'(x"cb"),u'(x"49"),u'(x"c3"),u'(x"06"),u'(x"85"),u'(x"df"),u'(x"00"),u'(x"cc"),u'(x"4f"),u'(x"df"),u'(x"cc"),
u'(x"04"),u'(x"df"),u'(x"c3"),u'(x"78"),u'(x"00"),u'(x"9f"),u'(x"cc"),u'(x"57"),u'(x"01"),u'(x"00"),u'(x"d7"),u'(x"cc"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"c4"),
u'(x"78"),u'(x"00"),u'(x"9f"),u'(x"cc"),u'(x"5f"),u'(x"7a"),u'(x"d7"),u'(x"cc"),u'(x"03"),u'(x"04"),u'(x"df"),u'(x"c5"),u'(x"78"),u'(x"00"),u'(x"9f"),u'(x"cc"),
u'(x"af"),u'(x"7f"),u'(x"02"),u'(x"00"),u'(x"6a"),u'(x"d7"),u'(x"cc"),u'(x"04"),u'(x"10"),u'(x"df"),u'(x"c6"),u'(x"78"),u'(x"00"),u'(x"d7"),u'(x"cc"),u'(x"02"),
u'(x"04"),u'(x"df"),u'(x"c7"),u'(x"78"),u'(x"00"),u'(x"9f"),u'(x"cc"),u'(x"77"),u'(x"ba"),u'(x"c6"),u'(x"fe"),u'(x"9f"),u'(x"ce"),u'(x"9f"),u'(x"d0"),u'(x"df"),
u'(x"02"),u'(x"d0"),u'(x"df"),u'(x"01"),u'(x"cc"),u'(x"c1"),u'(x"f2"),u'(x"04"),u'(x"44"),u'(x"09"),u'(x"df"),u'(x"02"),u'(x"cc"),u'(x"04"),u'(x"df"),u'(x"c8"),
u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"d0"),u'(x"06"),u'(x"97"),u'(x"aa"),u'(x"03"),u'(x"c4"),u'(x"2e"),u'(x"04"),u'(x"df"),u'(x"c9"),u'(x"78"),u'(x"00"),u'(x"9f"),
u'(x"cc"),u'(x"c6"),u'(x"ce"),u'(x"c1"),u'(x"f0"),u'(x"04"),u'(x"19"),u'(x"00"),u'(x"6e"),u'(x"df"),u'(x"01"),u'(x"cc"),u'(x"04"),u'(x"df"),u'(x"ca"),u'(x"78"),
u'(x"00"),u'(x"c6"),u'(x"d0"),u'(x"06"),u'(x"97"),u'(x"ff"),u'(x"03"),u'(x"c4"),u'(x"b4"),u'(x"04"),u'(x"df"),u'(x"cb"),u'(x"78"),u'(x"00"),u'(x"9f"),u'(x"cc"),
u'(x"c6"),u'(x"ce"),u'(x"c4"),u'(x"aa"),u'(x"c1"),u'(x"b4"),u'(x"11"),u'(x"df"),u'(x"04"),u'(x"cc"),u'(x"04"),u'(x"df"),u'(x"cc"),u'(x"78"),u'(x"00"),u'(x"c6"),
u'(x"d0"),u'(x"06"),u'(x"97"),u'(x"55"),u'(x"03"),u'(x"c4"),u'(x"ac"),u'(x"04"),u'(x"df"),u'(x"cd"),u'(x"78"),u'(x"00"),u'(x"9f"),u'(x"cc"),u'(x"c6"),u'(x"ce"),
u'(x"c4"),u'(x"ff"),u'(x"c1"),u'(x"6e"),u'(x"29"),u'(x"00"),u'(x"ec"),u'(x"df"),u'(x"03"),u'(x"cc"),u'(x"04"),u'(x"df"),u'(x"ce"),u'(x"78"),u'(x"00"),u'(x"c6"),
u'(x"d0"),u'(x"06"),u'(x"97"),u'(x"00"),u'(x"03"),u'(x"c4"),u'(x"ee"),u'(x"04"),u'(x"df"),u'(x"cf"),u'(x"78"),u'(x"00"),u'(x"9f"),u'(x"cc"),u'(x"c6"),u'(x"ce"),
u'(x"c4"),u'(x"55"),u'(x"c1"),u'(x"30"),u'(x"af"),u'(x"21"),u'(x"df"),u'(x"06"),u'(x"cc"),u'(x"04"),u'(x"df"),u'(x"d0"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"d0"),
u'(x"06"),u'(x"97"),u'(x"2e"),u'(x"03"),u'(x"c4"),u'(x"2a"),u'(x"04"),u'(x"df"),u'(x"d1"),u'(x"78"),u'(x"00"),u'(x"9f"),u'(x"cc"),u'(x"c6"),u'(x"ce"),u'(x"c4"),
u'(x"fb"),u'(x"c1"),u'(x"f2"),u'(x"39"),u'(x"f8"),u'(x"2a"),u'(x"df"),u'(x"05"),u'(x"cc"),u'(x"04"),u'(x"df"),u'(x"d2"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"d0"),
u'(x"06"),u'(x"97"),u'(x"ff"),u'(x"03"),u'(x"c4"),u'(x"6a"),u'(x"04"),u'(x"df"),u'(x"d3"),u'(x"78"),u'(x"00"),u'(x"9f"),u'(x"cc"),u'(x"c6"),u'(x"ce"),u'(x"c4"),
u'(x"2e"),u'(x"c1"),u'(x"b4"),u'(x"31"),u'(x"f8"),u'(x"df"),u'(x"07"),u'(x"cc"),u'(x"04"),u'(x"df"),u'(x"d4"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"d0"),u'(x"06"),
u'(x"97"),u'(x"fb"),u'(x"03"),u'(x"c4"),u'(x"ea"),u'(x"04"),u'(x"df"),u'(x"d5"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"ce"),u'(x"df"),u'(x"01"),u'(x"cc"),u'(x"9f"),
u'(x"ce"),u'(x"9f"),u'(x"d0"),u'(x"df"),u'(x"02"),u'(x"d0"),u'(x"c4"),u'(x"ff"),u'(x"17"),u'(x"a0"),u'(x"df"),u'(x"01"),u'(x"cc"),u'(x"09"),u'(x"c6"),u'(x"d0"),
u'(x"06"),u'(x"97"),u'(x"ff"),u'(x"03"),u'(x"17"),u'(x"74"),u'(x"04"),u'(x"df"),u'(x"d6"),u'(x"78"),u'(x"00"),u'(x"9f"),u'(x"cc"),u'(x"c4"),u'(x"55"),u'(x"c6"),
u'(x"ce"),u'(x"1f"),u'(x"de"),u'(x"00"),u'(x"d7"),u'(x"cc"),u'(x"03"),u'(x"09"),u'(x"c6"),u'(x"d0"),u'(x"06"),u'(x"97"),u'(x"55"),u'(x"03"),u'(x"17"),u'(x"10"),
u'(x"04"),u'(x"df"),u'(x"d7"),u'(x"78"),u'(x"00"),u'(x"9f"),u'(x"cc"),u'(x"c6"),u'(x"ce"),u'(x"c4"),u'(x"01"),u'(x"3f"),u'(x"02"),u'(x"00"),u'(x"10"),u'(x"d7"),
u'(x"cc"),u'(x"02"),u'(x"09"),u'(x"c6"),u'(x"d0"),u'(x"06"),u'(x"97"),u'(x"55"),u'(x"03"),u'(x"17"),u'(x"a6"),u'(x"04"),u'(x"df"),u'(x"d8"),u'(x"78"),u'(x"00"),
u'(x"9f"),u'(x"cc"),u'(x"c6"),u'(x"ce"),u'(x"c4"),u'(x"55"),u'(x"37"),u'(x"98"),u'(x"d7"),u'(x"cc"),u'(x"04"),u'(x"09"),u'(x"c6"),u'(x"d0"),u'(x"06"),u'(x"97"),
u'(x"01"),u'(x"03"),u'(x"17"),u'(x"da"),u'(x"04"),u'(x"df"),u'(x"d9"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"ce"),u'(x"c6"),u'(x"fe"),u'(x"e6"),u'(x"2e"),u'(x"c3"),
u'(x"4c"),u'(x"83"),u'(x"df"),u'(x"da"),u'(x"78"),u'(x"00"),u'(x"c3"),u'(x"2e"),u'(x"04"),u'(x"df"),u'(x"db"),u'(x"78"),u'(x"00"),u'(x"81"),u'(x"c5"),u'(x"6c"),
u'(x"46"),u'(x"86"),u'(x"df"),u'(x"dc"),u'(x"78"),u'(x"00"),u'(x"46"),u'(x"04"),u'(x"df"),u'(x"dd"),u'(x"78"),u'(x"00"),u'(x"46"),u'(x"df"),u'(x"00"),u'(x"fe"),
u'(x"c6"),u'(x"ff"),u'(x"c6"),u'(x"ff"),u'(x"04"),u'(x"df"),u'(x"de"),u'(x"78"),u'(x"00"),u'(x"06"),u'(x"c6"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"df"),u'(x"78"),
u'(x"00"),u'(x"c6"),u'(x"aa"),u'(x"c6"),u'(x"aa"),u'(x"04"),u'(x"df"),u'(x"e0"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"55"),u'(x"c6"),u'(x"55"),u'(x"04"),u'(x"df"),
u'(x"e1"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"c0"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"c6"),u'(x"ff"),u'(x"c6"),u'(x"ff"),u'(x"04"),u'(x"df"),u'(x"e2"),u'(x"78"),
u'(x"00"),u'(x"06"),u'(x"c6"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"e3"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"aa"),u'(x"c6"),u'(x"aa"),u'(x"04"),u'(x"df"),u'(x"e4"),
u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"55"),u'(x"c6"),u'(x"55"),u'(x"04"),u'(x"df"),u'(x"e5"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"80"),u'(x"1f"),u'(x"fe"),u'(x"c6"),
u'(x"fe"),u'(x"1f"),u'(x"c0"),u'(x"1f"),u'(x"80"),u'(x"1f"),u'(x"fe"),u'(x"f7"),u'(x"3e"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"c6"),u'(x"c0"),u'(x"04"),u'(x"df"),
u'(x"e6"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"c6"),u'(x"80"),u'(x"04"),u'(x"df"),u'(x"e7"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"fe"),u'(x"c6"),
u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"e8"),u'(x"78"),u'(x"00"),u'(x"77"),u'(x"bc"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"f7"),u'(x"36"),u'(x"ce"),u'(x"00"),u'(x"04"),
u'(x"df"),u'(x"e9"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"ce"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"ea"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"fe"),
u'(x"ce"),u'(x"32"),u'(x"04"),u'(x"df"),u'(x"eb"),u'(x"78"),u'(x"00"),u'(x"87"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"f7"),u'(x"36"),u'(x"ce"),u'(x"00"),u'(x"04"),
u'(x"df"),u'(x"ec"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"fe"),u'(x"ce"),u'(x"32"),u'(x"04"),u'(x"df"),u'(x"ed"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fe"),
u'(x"ce"),u'(x"7a"),u'(x"04"),u'(x"df"),u'(x"ee"),u'(x"78"),u'(x"00"),u'(x"87"),u'(x"ce"),u'(x"ba"),u'(x"04"),u'(x"df"),u'(x"ef"),u'(x"78"),u'(x"00"),u'(x"df"),
u'(x"00"),u'(x"fe"),u'(x"ce"),u'(x"7a"),u'(x"04"),u'(x"df"),u'(x"f0"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"fe"),u'(x"ce"),u'(x"32"),u'(x"04"),u'(x"df"),u'(x"f1"),
u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"87"),u'(x"bf"),u'(x"a4"),u'(x"c4"),u'(x"00"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"f2"),
u'(x"78"),u'(x"00"),u'(x"bf"),u'(x"a9"),u'(x"c4"),u'(x"00"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"f3"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"44"),
u'(x"bf"),u'(x"a4"),u'(x"c4"),u'(x"00"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"f4"),u'(x"78"),u'(x"00"),u'(x"bf"),u'(x"a9"),u'(x"c4"),u'(x"00"),
u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"f5"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"44"),u'(x"bf"),u'(x"a4"),u'(x"c4"),u'(x"ff"),u'(x"03"),u'(x"02"),
u'(x"01"),u'(x"04"),u'(x"df"),u'(x"f6"),u'(x"78"),u'(x"00"),u'(x"44"),u'(x"bf"),u'(x"a9"),u'(x"c4"),u'(x"ff"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),
u'(x"f7"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"bf"),u'(x"a6"),u'(x"c4"),u'(x"00"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"f8"),u'(x"78"),u'(x"00"),
u'(x"bf"),u'(x"a1"),u'(x"c4"),u'(x"37"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"f9"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"ff"),u'(x"af"),u'(x"b1"),
u'(x"84"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"fa"),u'(x"78"),u'(x"00"),u'(x"af"),u'(x"84"),u'(x"0b"),u'(x"0a"),u'(x"c4"),u'(x"08"),u'(x"07"),
u'(x"bf"),u'(x"aa"),u'(x"c4"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"fb"),u'(x"78"),u'(x"00"),u'(x"bf"),u'(x"a4"),u'(x"04"),u'(x"03"),u'(x"02"),
u'(x"01"),u'(x"04"),u'(x"df"),u'(x"fc"),u'(x"78"),u'(x"00"),u'(x"44"),u'(x"bf"),u'(x"c4"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"fd"),u'(x"78"),
u'(x"00"),u'(x"bf"),u'(x"c4"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"fe"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"ff"),u'(x"c1"),u'(x"01"),u'(x"af"),u'(x"01"),
u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"ff"),u'(x"78"),u'(x"00"),u'(x"84"),u'(x"01"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"00"),u'(x"78"),
u'(x"00"),u'(x"01"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"01"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"ff"),u'(x"bf"),u'(x"44"),u'(x"03"),u'(x"02"),u'(x"01"),
u'(x"04"),u'(x"df"),u'(x"02"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"ff"),u'(x"bf"),u'(x"a2"),u'(x"44"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"03"),
u'(x"78"),u'(x"00"),u'(x"bf"),u'(x"44"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"04"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"ff"),u'(x"af"),u'(x"04"),u'(x"03"),
u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"05"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"af"),u'(x"04"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"06"),
u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"ff"),u'(x"c1"),u'(x"00"),u'(x"af"),u'(x"01"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"07"),u'(x"78"),u'(x"00"),
u'(x"af"),u'(x"41"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"08"),u'(x"78"),u'(x"00"),u'(x"bf"),u'(x"41"),u'(x"04"),u'(x"df"),u'(x"09"),u'(x"78"),
u'(x"00"),u'(x"c4"),u'(x"fd"),u'(x"af"),u'(x"c4"),u'(x"ef"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"0a"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"05"),
u'(x"af"),u'(x"c4"),u'(x"0a"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"0b"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"00"),u'(x"af"),u'(x"84"),u'(x"06"),
u'(x"05"),u'(x"b1"),u'(x"84"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"0c"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"bf"),u'(x"a1"),u'(x"84"),u'(x"08"),u'(x"07"),
u'(x"06"),u'(x"b1"),u'(x"84"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"0d"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"00"),u'(x"af"),u'(x"44"),u'(x"02"),
u'(x"01"),u'(x"04"),u'(x"df"),u'(x"0e"),u'(x"78"),u'(x"00"),u'(x"44"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"0f"),u'(x"78"),u'(x"00"),u'(x"44"),u'(x"03"),
u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"10"),u'(x"78"),u'(x"00"),u'(x"44"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"11"),u'(x"78"),u'(x"00"),u'(x"c4"),
u'(x"03"),u'(x"af"),u'(x"04"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"12"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"13"),
u'(x"78"),u'(x"00"),u'(x"04"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"14"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"15"),
u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"55"),u'(x"a1"),u'(x"01"),u'(x"01"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"16"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"aa"),u'(x"04"),
u'(x"df"),u'(x"17"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"aa"),u'(x"a1"),u'(x"41"),u'(x"41"),u'(x"41"),u'(x"04"),u'(x"df"),u'(x"18"),u'(x"78"),u'(x"00"),u'(x"c1"),
u'(x"52"),u'(x"04"),u'(x"df"),u'(x"19"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"00"),u'(x"af"),u'(x"c4"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"1a"),u'(x"78"),
u'(x"00"),u'(x"c4"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"1b"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"1c"),
u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"1d"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"e1"),u'(x"af"),u'(x"84"),u'(x"02"),u'(x"01"),
u'(x"04"),u'(x"df"),u'(x"1e"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"01"),u'(x"84"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"1f"),u'(x"78"),u'(x"00"),u'(x"84"),
u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"20"),u'(x"78"),u'(x"00"),u'(x"84"),u'(x"05"),u'(x"04"),u'(x"03"),u'(x"c4"),u'(x"0e"),u'(x"04"),u'(x"df"),u'(x"21"),
u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"2e"),u'(x"01"),u'(x"af"),u'(x"c4"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"22"),u'(x"78"),u'(x"00"),u'(x"44"),
u'(x"bf"),u'(x"c4"),u'(x"05"),u'(x"04"),u'(x"03"),u'(x"02"),u'(x"44"),u'(x"04"),u'(x"df"),u'(x"23"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"2e"),u'(x"c1"),u'(x"55"),
u'(x"af"),u'(x"44"),u'(x"03"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"24"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"aa"),u'(x"bf"),u'(x"44"),u'(x"03"),u'(x"02"),
u'(x"01"),u'(x"04"),u'(x"df"),u'(x"25"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"06"),u'(x"05"),u'(x"04"),u'(x"03"),u'(x"c4"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"26"),
u'(x"78"),u'(x"00"),u'(x"04"),u'(x"af"),u'(x"b9"),u'(x"c4"),u'(x"05"),u'(x"04"),u'(x"03"),u'(x"02"),u'(x"84"),u'(x"04"),u'(x"df"),u'(x"27"),u'(x"78"),u'(x"00"),
u'(x"bf"),u'(x"a8"),u'(x"04"),u'(x"cc"),u'(x"2d"),u'(x"cc"),u'(x"05"),u'(x"04"),u'(x"03"),u'(x"02"),u'(x"cc"),u'(x"04"),u'(x"df"),u'(x"28"),u'(x"78"),u'(x"00"),
u'(x"c0"),u'(x"ff"),u'(x"04"),u'(x"c0"),u'(x"c0"),u'(x"04"),u'(x"df"),u'(x"29"),u'(x"78"),u'(x"00"),u'(x"00"),u'(x"c0"),u'(x"ff"),u'(x"c0"),u'(x"c0"),u'(x"ff"),
u'(x"04"),u'(x"df"),u'(x"2a"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"a3"),u'(x"c4"),u'(x"db"),u'(x"bf"),u'(x"01"),u'(x"06"),u'(x"05"),u'(x"04"),u'(x"03"),u'(x"57"),
u'(x"78"),u'(x"04"),u'(x"df"),u'(x"2b"),u'(x"78"),u'(x"00"),u'(x"42"),u'(x"af"),u'(x"02"),u'(x"05"),u'(x"04"),u'(x"03"),u'(x"97"),u'(x"a3"),u'(x"04"),u'(x"df"),
u'(x"2c"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"6d"),u'(x"bf"),u'(x"10"),u'(x"0f"),u'(x"0e"),u'(x"0d"),u'(x"05"),u'(x"05"),u'(x"04"),u'(x"03"),u'(x"02"),u'(x"77"),
u'(x"14"),u'(x"df"),u'(x"2d"),u'(x"78"),u'(x"00"),u'(x"77"),u'(x"08"),u'(x"df"),u'(x"2e"),u'(x"78"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"2f"),
u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"be"),u'(x"df"),u'(x"aa"),u'(x"fc"),u'(x"c5"),u'(x"c2"),u'(x"e6"),u'(x"1f"),u'(x"bf"),u'(x"4e"),u'(x"df"),u'(x"30"),u'(x"78"),
u'(x"00"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"31"),u'(x"78"),u'(x"00"),u'(x"c5"),u'(x"aa"),u'(x"04"),u'(x"df"),u'(x"32"),u'(x"78"),u'(x"00"),u'(x"97"),
u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"33"),u'(x"78"),u'(x"00"),u'(x"e6"),u'(x"55"),u'(x"e6"),u'(x"00"),u'(x"85"),u'(x"f7"),u'(x"04"),u'(x"77"),u'(x"0c"),u'(x"af"),
u'(x"85"),u'(x"df"),u'(x"34"),u'(x"78"),u'(x"00"),u'(x"02"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"35"),u'(x"78"),u'(x"00"),u'(x"97"),u'(x"fe"),u'(x"04"),u'(x"df"),
u'(x"36"),u'(x"78"),u'(x"00"),u'(x"c5"),u'(x"55"),u'(x"04"),u'(x"df"),u'(x"37"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"0f"),u'(x"fe"),u'(x"af"),u'(x"df"),u'(x"00"),
u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"38"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"0f"),u'(x"fe"),u'(x"a1"),u'(x"df"),u'(x"0e"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"39"),
u'(x"78"),u'(x"00"),u'(x"df"),u'(x"0f"),u'(x"fe"),u'(x"a8"),u'(x"df"),u'(x"07"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"3a"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"0f"),
u'(x"fe"),u'(x"a2"),u'(x"df"),u'(x"0d"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"3b"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"0f"),u'(x"fe"),u'(x"a4"),u'(x"df"),u'(x"0b"),
u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"3c"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"bf"),u'(x"df"),u'(x"0f"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"3d"),
u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"b1"),u'(x"df"),u'(x"01"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"3e"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),
u'(x"fe"),u'(x"b8"),u'(x"df"),u'(x"08"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"3f"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"b2"),u'(x"df"),u'(x"02"),
u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"40"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"b4"),u'(x"df"),u'(x"04"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"41"),
u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"bf"),u'(x"a3"),u'(x"df"),u'(x"0c"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"42"),u'(x"78"),u'(x"00"),u'(x"bf"),
u'(x"a5"),u'(x"df"),u'(x"0a"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"43"),u'(x"78"),u'(x"00"),u'(x"bf"),u'(x"a6"),u'(x"df"),u'(x"09"),u'(x"fe"),u'(x"04"),u'(x"df"),
u'(x"44"),u'(x"78"),u'(x"00"),u'(x"bf"),u'(x"a7"),u'(x"df"),u'(x"08"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"45"),u'(x"78"),u'(x"00"),u'(x"bf"),u'(x"a9"),u'(x"df"),
u'(x"06"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"46"),u'(x"78"),u'(x"00"),u'(x"bf"),u'(x"aa"),u'(x"df"),u'(x"05"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"47"),u'(x"78"),
u'(x"00"),u'(x"bf"),u'(x"ab"),u'(x"df"),u'(x"04"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"48"),u'(x"78"),u'(x"00"),u'(x"bf"),u'(x"ac"),u'(x"df"),u'(x"03"),u'(x"fe"),
u'(x"04"),u'(x"df"),u'(x"49"),u'(x"78"),u'(x"00"),u'(x"bf"),u'(x"ad"),u'(x"df"),u'(x"02"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"4a"),u'(x"78"),u'(x"00"),u'(x"bf"),
u'(x"ae"),u'(x"df"),u'(x"01"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"4b"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"b3"),u'(x"df"),u'(x"03"),u'(x"fe"),
u'(x"04"),u'(x"df"),u'(x"4c"),u'(x"78"),u'(x"00"),u'(x"af"),u'(x"b5"),u'(x"df"),u'(x"05"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"4d"),u'(x"78"),u'(x"00"),u'(x"af"),
u'(x"b6"),u'(x"df"),u'(x"06"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"4e"),u'(x"78"),u'(x"00"),u'(x"af"),u'(x"b7"),u'(x"df"),u'(x"07"),u'(x"fe"),u'(x"04"),u'(x"df"),
u'(x"4f"),u'(x"78"),u'(x"00"),u'(x"af"),u'(x"b9"),u'(x"df"),u'(x"09"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"50"),u'(x"78"),u'(x"00"),u'(x"af"),u'(x"ba"),u'(x"df"),
u'(x"0a"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"51"),u'(x"78"),u'(x"00"),u'(x"af"),u'(x"bb"),u'(x"df"),u'(x"0b"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"52"),u'(x"78"),
u'(x"00"),u'(x"af"),u'(x"bc"),u'(x"df"),u'(x"0c"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"53"),u'(x"78"),u'(x"00"),u'(x"af"),u'(x"bd"),u'(x"df"),u'(x"0d"),u'(x"fe"),
u'(x"04"),u'(x"df"),u'(x"54"),u'(x"78"),u'(x"00"),u'(x"af"),u'(x"be"),u'(x"df"),u'(x"0e"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"55"),u'(x"78"),u'(x"00"),u'(x"af"),
u'(x"04"),u'(x"df"),u'(x"56"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"57"),u'(x"78"),u'(x"00"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"58"),u'(x"78"),u'(x"00"),
u'(x"01"),u'(x"04"),u'(x"df"),u'(x"59"),u'(x"78"),u'(x"00"),u'(x"b4"),u'(x"04"),u'(x"df"),u'(x"5a"),u'(x"78"),u'(x"00"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"5b"),
u'(x"78"),u'(x"00"),u'(x"af"),u'(x"b8"),u'(x"04"),u'(x"df"),u'(x"5c"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"5d"),u'(x"78"),u'(x"00"),u'(x"01"),u'(x"04"),
u'(x"df"),u'(x"5e"),u'(x"78"),u'(x"00"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"5f"),u'(x"78"),u'(x"00"),u'(x"af"),u'(x"b2"),u'(x"04"),u'(x"df"),u'(x"60"),u'(x"78"),
u'(x"00"),u'(x"04"),u'(x"df"),u'(x"61"),u'(x"78"),u'(x"00"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"62"),u'(x"78"),u'(x"00"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"63"),
u'(x"78"),u'(x"00"),u'(x"af"),u'(x"ba"),u'(x"04"),u'(x"df"),u'(x"64"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"65"),u'(x"78"),u'(x"00"),u'(x"01"),u'(x"04"),
u'(x"df"),u'(x"66"),u'(x"78"),u'(x"00"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"67"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"c0"),u'(x"01"),u'(x"c1"),
u'(x"02"),u'(x"c2"),u'(x"03"),u'(x"c3"),u'(x"04"),u'(x"c4"),u'(x"05"),u'(x"c5"),u'(x"06"),u'(x"9f"),u'(x"c4"),u'(x"df"),u'(x"0f"),u'(x"ca"),u'(x"bf"),u'(x"a0"),
u'(x"a0"),u'(x"a0"),u'(x"f7"),u'(x"32"),u'(x"9f"),u'(x"c4"),u'(x"04"),u'(x"df"),u'(x"68"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"ca"),u'(x"af"),u'(x"b0"),
u'(x"b0"),u'(x"b0"),u'(x"f7"),u'(x"12"),u'(x"9f"),u'(x"c4"),u'(x"04"),u'(x"df"),u'(x"69"),u'(x"78"),u'(x"00"),u'(x"77"),u'(x"66"),u'(x"df"),u'(x"ca"),u'(x"fe"),
u'(x"04"),u'(x"df"),u'(x"6a"),u'(x"78"),u'(x"00"),u'(x"c0"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"6b"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"02"),u'(x"04"),u'(x"df"),
u'(x"6c"),u'(x"78"),u'(x"00"),u'(x"c2"),u'(x"03"),u'(x"04"),u'(x"df"),u'(x"6d"),u'(x"78"),u'(x"00"),u'(x"c3"),u'(x"04"),u'(x"04"),u'(x"df"),u'(x"6e"),u'(x"78"),
u'(x"00"),u'(x"c4"),u'(x"05"),u'(x"04"),u'(x"df"),u'(x"6f"),u'(x"78"),u'(x"00"),u'(x"c5"),u'(x"06"),u'(x"04"),u'(x"df"),u'(x"70"),u'(x"78"),u'(x"00"),u'(x"87"),
u'(x"00"),u'(x"01"),u'(x"02"),u'(x"03"),u'(x"04"),u'(x"05"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"71"),u'(x"78"),
u'(x"00"),u'(x"c0"),u'(x"ff"),u'(x"01"),u'(x"42"),u'(x"83"),u'(x"c4"),u'(x"05"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"04"),u'(x"df"),
u'(x"72"),u'(x"78"),u'(x"00"),u'(x"c0"),u'(x"04"),u'(x"df"),u'(x"73"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"04"),u'(x"df"),u'(x"74"),u'(x"78"),u'(x"00"),u'(x"c2"),
u'(x"04"),u'(x"df"),u'(x"75"),u'(x"78"),u'(x"00"),u'(x"c3"),u'(x"04"),u'(x"df"),u'(x"76"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"04"),u'(x"df"),u'(x"77"),u'(x"78"),
u'(x"00"),u'(x"c5"),u'(x"04"),u'(x"df"),u'(x"78"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"00"),u'(x"01"),u'(x"02"),u'(x"03"),u'(x"04"),u'(x"05"),
u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"c0"),u'(x"ff"),u'(x"01"),u'(x"42"),u'(x"83"),u'(x"c4"),u'(x"05"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"c0"),u'(x"04"),u'(x"df"),
u'(x"79"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"04"),u'(x"df"),u'(x"7a"),u'(x"78"),u'(x"00"),u'(x"c2"),u'(x"04"),u'(x"df"),u'(x"7b"),u'(x"78"),u'(x"00"),u'(x"c3"),
u'(x"04"),u'(x"df"),u'(x"7c"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"04"),u'(x"df"),u'(x"7d"),u'(x"78"),u'(x"00"),u'(x"c5"),u'(x"04"),u'(x"df"),u'(x"7e"),u'(x"78"),
u'(x"00"),u'(x"c0"),u'(x"ff"),u'(x"17"),u'(x"ff"),u'(x"04"),u'(x"df"),u'(x"7f"),u'(x"78"),u'(x"00"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"80"),
u'(x"78"),u'(x"00"),u'(x"c0"),u'(x"aa"),u'(x"17"),u'(x"aa"),u'(x"04"),u'(x"df"),u'(x"81"),u'(x"78"),u'(x"00"),u'(x"c0"),u'(x"55"),u'(x"17"),u'(x"55"),u'(x"04"),
u'(x"df"),u'(x"82"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"ff"),u'(x"57"),u'(x"ff"),u'(x"04"),u'(x"df"),u'(x"83"),u'(x"78"),u'(x"00"),u'(x"01"),u'(x"57"),u'(x"00"),
u'(x"04"),u'(x"df"),u'(x"84"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"aa"),u'(x"57"),u'(x"aa"),u'(x"04"),u'(x"df"),u'(x"85"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"55"),
u'(x"57"),u'(x"55"),u'(x"04"),u'(x"df"),u'(x"86"),u'(x"78"),u'(x"00"),u'(x"c2"),u'(x"ff"),u'(x"97"),u'(x"ff"),u'(x"04"),u'(x"df"),u'(x"87"),u'(x"78"),u'(x"00"),
u'(x"02"),u'(x"97"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"88"),u'(x"78"),u'(x"00"),u'(x"c2"),u'(x"aa"),u'(x"97"),u'(x"aa"),u'(x"04"),u'(x"df"),u'(x"89"),u'(x"78"),
u'(x"00"),u'(x"c2"),u'(x"55"),u'(x"97"),u'(x"55"),u'(x"04"),u'(x"df"),u'(x"8a"),u'(x"78"),u'(x"00"),u'(x"c3"),u'(x"ff"),u'(x"d7"),u'(x"ff"),u'(x"04"),u'(x"df"),
u'(x"8b"),u'(x"78"),u'(x"00"),u'(x"03"),u'(x"d7"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"8c"),u'(x"78"),u'(x"00"),u'(x"c3"),u'(x"aa"),u'(x"d7"),u'(x"aa"),u'(x"04"),
u'(x"df"),u'(x"8d"),u'(x"78"),u'(x"00"),u'(x"c3"),u'(x"55"),u'(x"d7"),u'(x"55"),u'(x"04"),u'(x"df"),u'(x"8e"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"ff"),u'(x"17"),
u'(x"ff"),u'(x"04"),u'(x"df"),u'(x"8f"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"17"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"90"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"aa"),
u'(x"17"),u'(x"aa"),u'(x"04"),u'(x"df"),u'(x"91"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"55"),u'(x"17"),u'(x"55"),u'(x"04"),u'(x"df"),u'(x"92"),u'(x"78"),u'(x"00"),
u'(x"c5"),u'(x"ff"),u'(x"57"),u'(x"ff"),u'(x"04"),u'(x"df"),u'(x"93"),u'(x"78"),u'(x"00"),u'(x"05"),u'(x"57"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"94"),u'(x"78"),
u'(x"00"),u'(x"c5"),u'(x"aa"),u'(x"57"),u'(x"aa"),u'(x"04"),u'(x"df"),u'(x"95"),u'(x"78"),u'(x"00"),u'(x"c5"),u'(x"55"),u'(x"57"),u'(x"55"),u'(x"04"),u'(x"df"),
u'(x"96"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"04"),u'(x"c1"),u'(x"be"),u'(x"c2"),u'(x"c6"),u'(x"c3"),u'(x"cc"),u'(x"5f"),u'(x"fe"),u'(x"c4"),
u'(x"d2"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"97"),u'(x"78"),u'(x"00"),u'(x"13"),u'(x"04"),u'(x"df"),u'(x"98"),u'(x"78"),u'(x"00"),u'(x"57"),u'(x"ff"),u'(x"ed"),
u'(x"c1"),u'(x"be"),u'(x"c2"),u'(x"c6"),u'(x"c3"),u'(x"cc"),u'(x"85"),u'(x"5f"),u'(x"fe"),u'(x"c6"),u'(x"ca"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"99"),u'(x"78"),
u'(x"00"),u'(x"8b"),u'(x"04"),u'(x"df"),u'(x"9a"),u'(x"78"),u'(x"00"),u'(x"46"),u'(x"c1"),u'(x"be"),u'(x"c2"),u'(x"c6"),u'(x"c3"),u'(x"d2"),u'(x"1f"),u'(x"ca"),
u'(x"c4"),u'(x"ca"),u'(x"5f"),u'(x"fe"),u'(x"d4"),u'(x"d2"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"9b"),u'(x"78"),u'(x"00"),u'(x"17"),u'(x"cb"),u'(x"04"),u'(x"df"),
u'(x"9c"),u'(x"78"),u'(x"00"),u'(x"d3"),u'(x"ca"),u'(x"04"),u'(x"df"),u'(x"9d"),u'(x"78"),u'(x"00"),u'(x"57"),u'(x"ff"),u'(x"e3"),u'(x"77"),u'(x"1a"),u'(x"87"),
u'(x"00"),u'(x"2f"),u'(x"ff"),u'(x"89"),u'(x"04"),u'(x"21"),u'(x"87"),u'(x"00"),u'(x"2f"),u'(x"87"),u'(x"00"),u'(x"2f"),u'(x"a0"),u'(x"df"),u'(x"00"),u'(x"fe"),
u'(x"c1"),u'(x"b8"),u'(x"c2"),u'(x"a8"),u'(x"43"),u'(x"f7"),u'(x"5e"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"c6"),u'(x"80"),u'(x"c1"),u'(x"b8"),u'(x"c2"),u'(x"b0"),
u'(x"43"),u'(x"f7"),u'(x"46"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"c1"),u'(x"a4"),u'(x"c2"),u'(x"b0"),u'(x"c3"),u'(x"b8"),u'(x"44"),u'(x"f7"),u'(x"54"),u'(x"df"),
u'(x"00"),u'(x"fe"),u'(x"c1"),u'(x"a4"),u'(x"c2"),u'(x"a8"),u'(x"c3"),u'(x"b8"),u'(x"1f"),u'(x"fe"),u'(x"17"),u'(x"0a"),u'(x"df"),u'(x"0a"),u'(x"fe"),u'(x"04"),
u'(x"df"),u'(x"9e"),u'(x"78"),u'(x"00"),u'(x"77"),u'(x"74"),u'(x"45"),u'(x"05"),u'(x"d2"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"9f"),u'(x"78"),u'(x"00"),u'(x"c5"),
u'(x"04"),u'(x"df"),u'(x"a0"),u'(x"78"),u'(x"00"),u'(x"97"),u'(x"ff"),u'(x"ee"),u'(x"87"),u'(x"11"),u'(x"d2"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"a1"),u'(x"78"),
u'(x"00"),u'(x"13"),u'(x"04"),u'(x"df"),u'(x"a2"),u'(x"78"),u'(x"00"),u'(x"44"),u'(x"04"),u'(x"df"),u'(x"a3"),u'(x"78"),u'(x"00"),u'(x"83"),u'(x"97"),u'(x"ff"),
u'(x"e8"),u'(x"87"),u'(x"ff"),u'(x"aa"),u'(x"ef"),u'(x"00"),u'(x"aa"),u'(x"ff"),u'(x"0f"),u'(x"00"),u'(x"0a"),u'(x"05"),u'(x"ff"),u'(x"00"),u'(x"aa"),u'(x"55"),
u'(x"77"),u'(x"6a"),u'(x"e6"),u'(x"08"),u'(x"df"),u'(x"26"),u'(x"08"),u'(x"c0"),u'(x"ff"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"07"),u'(x"df"),u'(x"00"),u'(x"fe"),
u'(x"04"),u'(x"df"),u'(x"a4"),u'(x"78"),u'(x"00"),u'(x"17"),u'(x"49"),u'(x"04"),u'(x"df"),u'(x"a5"),u'(x"78"),u'(x"00"),u'(x"c0"),u'(x"ff"),u'(x"bf"),u'(x"07"),
u'(x"df"),u'(x"0f"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"a6"),u'(x"78"),u'(x"00"),u'(x"17"),u'(x"49"),u'(x"04"),u'(x"df"),u'(x"a7"),u'(x"78"),u'(x"00"),u'(x"9f"),
u'(x"08"),u'(x"77"),u'(x"08"),u'(x"df"),u'(x"a8"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"f6"),u'(x"1f"),u'(x"fe"),u'(x"e6"),u'(x"04"),u'(x"e6"),u'(x"06"),u'(x"e6"),
u'(x"08"),u'(x"e6"),u'(x"0a"),u'(x"df"),u'(x"72"),u'(x"04"),u'(x"1f"),u'(x"06"),u'(x"df"),u'(x"72"),u'(x"08"),u'(x"1f"),u'(x"0a"),u'(x"df"),u'(x"00"),u'(x"fe"),
u'(x"c6"),u'(x"80"),u'(x"00"),u'(x"df"),u'(x"a9"),u'(x"78"),u'(x"00"),u'(x"77"),u'(x"3e"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"aa"),u'(x"78"),
u'(x"00"),u'(x"df"),u'(x"80"),u'(x"f6"),u'(x"05"),u'(x"04"),u'(x"df"),u'(x"ab"),u'(x"78"),u'(x"00"),u'(x"97"),u'(x"66"),u'(x"04"),u'(x"df"),u'(x"ac"),u'(x"78"),
u'(x"00"),u'(x"97"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"ad"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"f6"),u'(x"9f"),u'(x"0a"),u'(x"9f"),u'(x"08"),u'(x"9f"),u'(x"06"),
u'(x"9f"),u'(x"04"),u'(x"df"),u'(x"e0"),u'(x"fe"),u'(x"df"),u'(x"00"),u'(x"7a"),u'(x"df"),u'(x"3f"),u'(x"4e"),u'(x"1f"),u'(x"fa"),u'(x"d7"),u'(x"fa"),u'(x"00"),
u'(x"04"),u'(x"df"),u'(x"ae"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fa"),u'(x"df"),u'(x"aa"),u'(x"fa"),u'(x"04"),u'(x"df"),u'(x"af"),u'(x"78"),u'(x"00"),
u'(x"df"),u'(x"00"),u'(x"fa"),u'(x"df"),u'(x"cc"),u'(x"fa"),u'(x"04"),u'(x"df"),u'(x"b0"),u'(x"78"),u'(x"00"),u'(x"bf"),u'(x"05"),u'(x"df"),u'(x"ef"),u'(x"fe"),
u'(x"04"),u'(x"df"),u'(x"b1"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"7a"),u'(x"c1"),u'(x"7e"),u'(x"c1"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"b2"),u'(x"78"),u'(x"00"),
u'(x"df"),u'(x"00"),u'(x"4e"),u'(x"04"),u'(x"df"),u'(x"b3"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fa"),u'(x"04"),u'(x"df"),u'(x"b4"),u'(x"78"),u'(x"00"),
u'(x"c2"),u'(x"04"),u'(x"c3"),u'(x"06"),u'(x"c4"),u'(x"08"),u'(x"c5"),u'(x"0a"),u'(x"df"),u'(x"f0"),u'(x"04"),u'(x"df"),u'(x"e0"),u'(x"06"),u'(x"df"),u'(x"f0"),
u'(x"08"),u'(x"df"),u'(x"e0"),u'(x"0a"),u'(x"df"),u'(x"e0"),u'(x"fe"),u'(x"df"),u'(x"00"),u'(x"7a"),u'(x"df"),u'(x"3f"),u'(x"4e"),u'(x"df"),u'(x"00"),u'(x"fa"),
u'(x"bf"),u'(x"05"),u'(x"df"),u'(x"ef"),u'(x"fe"),u'(x"05"),u'(x"00"),u'(x"df"),u'(x"b5"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"7a"),u'(x"c1"),u'(x"7e"),u'(x"c1"),
u'(x"00"),u'(x"05"),u'(x"00"),u'(x"df"),u'(x"b6"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"0f"),u'(x"4e"),u'(x"05"),u'(x"00"),u'(x"df"),u'(x"b7"),u'(x"78"),u'(x"00"),
u'(x"df"),u'(x"cc"),u'(x"fa"),u'(x"05"),u'(x"df"),u'(x"b8"),u'(x"78"),u'(x"00"),u'(x"02"),u'(x"1f"),u'(x"fa"),u'(x"1f"),u'(x"fe"),u'(x"9f"),u'(x"04"),u'(x"df"),
u'(x"06"),u'(x"1f"),u'(x"08"),u'(x"5f"),u'(x"0a"),u'(x"c5"),u'(x"08"),u'(x"c1"),u'(x"ae"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"f7"),u'(x"38"),u'(x"5f"),u'(x"fe"),
u'(x"04"),u'(x"df"),u'(x"b9"),u'(x"78"),u'(x"00"),u'(x"4d"),u'(x"c5"),u'(x"08"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"c6"),u'(x"80"),u'(x"f7"),u'(x"16"),u'(x"df"),
u'(x"0f"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"ba"),u'(x"78"),u'(x"00"),u'(x"50"),u'(x"77"),u'(x"6a"),u'(x"57"),u'(x"08"),u'(x"03"),u'(x"bf"),u'(x"98"),u'(x"26"),
u'(x"57"),u'(x"07"),u'(x"03"),u'(x"bf"),u'(x"99"),u'(x"20"),u'(x"57"),u'(x"06"),u'(x"03"),u'(x"bf"),u'(x"9a"),u'(x"1a"),u'(x"57"),u'(x"05"),u'(x"03"),u'(x"bf"),
u'(x"9b"),u'(x"14"),u'(x"57"),u'(x"04"),u'(x"03"),u'(x"bf"),u'(x"9c"),u'(x"0e"),u'(x"57"),u'(x"03"),u'(x"03"),u'(x"bf"),u'(x"9d"),u'(x"08"),u'(x"57"),u'(x"02"),
u'(x"03"),u'(x"bf"),u'(x"9e"),u'(x"02"),u'(x"bf"),u'(x"9f"),u'(x"87"),u'(x"0f"),u'(x"2f"),u'(x"4f"),u'(x"6f"),u'(x"8f"),u'(x"af"),u'(x"cf"),u'(x"ef"),u'(x"1f"),
u'(x"fe"),u'(x"c3"),u'(x"0a"),u'(x"c1"),u'(x"00"),u'(x"c0"),u'(x"4e"),u'(x"11"),u'(x"c2"),u'(x"e6"),u'(x"08"),u'(x"df"),u'(x"62"),u'(x"08"),u'(x"00"),u'(x"c1"),
u'(x"00"),u'(x"c2"),u'(x"08"),u'(x"c3"),u'(x"0e"),u'(x"44"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"b2"),u'(x"91"),u'(x"9f"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"bb"),
u'(x"78"),u'(x"00"),u'(x"0b"),u'(x"04"),u'(x"df"),u'(x"bc"),u'(x"78"),u'(x"00"),u'(x"84"),u'(x"84"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"bd"),u'(x"78"),u'(x"00"),
u'(x"cb"),u'(x"01"),u'(x"e1"),u'(x"04"),u'(x"df"),u'(x"be"),u'(x"78"),u'(x"00"),u'(x"81"),u'(x"81"),u'(x"57"),u'(x"ff"),u'(x"d9"),u'(x"df"),u'(x"6a"),u'(x"08"),
u'(x"81"),u'(x"df"),u'(x"bf"),u'(x"78"),u'(x"00"),u'(x"77"),u'(x"20"),u'(x"84"),u'(x"00"),u'(x"01"),u'(x"ff"),u'(x"08"),u'(x"04"),u'(x"01"),u'(x"84"),u'(x"00"),
u'(x"01"),u'(x"df"),u'(x"c0"),u'(x"78"),u'(x"00"),u'(x"d6"),u'(x"d6"),u'(x"9f"),u'(x"08"),u'(x"1f"),u'(x"fe"),u'(x"c3"),u'(x"0a"),u'(x"c1"),u'(x"00"),u'(x"c0"),
u'(x"0c"),u'(x"11"),u'(x"c2"),u'(x"e6"),u'(x"08"),u'(x"df"),u'(x"20"),u'(x"08"),u'(x"c1"),u'(x"00"),u'(x"c2"),u'(x"08"),u'(x"c3"),u'(x"0e"),u'(x"84"),u'(x"df"),
u'(x"00"),u'(x"fe"),u'(x"40"),u'(x"d7"),u'(x"0e"),u'(x"01"),u'(x"02"),u'(x"b1"),u'(x"01"),u'(x"a1"),u'(x"b2"),u'(x"d2"),u'(x"df"),u'(x"fe"),u'(x"04"),u'(x"df"),
u'(x"c1"),u'(x"78"),u'(x"00"),u'(x"40"),u'(x"04"),u'(x"df"),u'(x"c2"),u'(x"78"),u'(x"00"),u'(x"84"),u'(x"84"),u'(x"84"),u'(x"04"),u'(x"df"),u'(x"c3"),u'(x"78"),
u'(x"00"),u'(x"62"),u'(x"04"),u'(x"df"),u'(x"c4"),u'(x"78"),u'(x"00"),u'(x"82"),u'(x"82"),u'(x"57"),u'(x"ff"),u'(x"d3"),u'(x"df"),u'(x"28"),u'(x"08"),u'(x"c2"),
u'(x"df"),u'(x"c5"),u'(x"78"),u'(x"00"),u'(x"77"),u'(x"20"),u'(x"84"),u'(x"00"),u'(x"01"),u'(x"ff"),u'(x"ff"),u'(x"ff"),u'(x"ff"),u'(x"09"),u'(x"04"),u'(x"00"),
u'(x"df"),u'(x"c6"),u'(x"78"),u'(x"00"),u'(x"d6"),u'(x"d6"),u'(x"9f"),u'(x"08"),u'(x"1f"),u'(x"fe"),u'(x"c1"),u'(x"06"),u'(x"5f"),u'(x"ca"),u'(x"df"),u'(x"02"),
u'(x"ca"),u'(x"c3"),u'(x"92"),u'(x"42"),u'(x"bf"),u'(x"b1"),u'(x"02"),u'(x"5f"),u'(x"04"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"c7"),u'(x"78"),u'(x"00"),u'(x"43"),
u'(x"06"),u'(x"04"),u'(x"df"),u'(x"c8"),u'(x"78"),u'(x"00"),u'(x"42"),u'(x"08"),u'(x"04"),u'(x"df"),u'(x"c9"),u'(x"78"),u'(x"00"),u'(x"7f"),u'(x"02"),u'(x"4a"),
u'(x"04"),u'(x"df"),u'(x"ca"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"0a"),u'(x"57"),u'(x"9c"),u'(x"d2"),u'(x"c1"),u'(x"06"),u'(x"42"),u'(x"c6"),u'(x"fe"),u'(x"c4"),
u'(x"04"),u'(x"45"),u'(x"bf"),u'(x"71"),u'(x"02"),u'(x"5f"),u'(x"04"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"cb"),u'(x"78"),u'(x"00"),u'(x"45"),u'(x"06"),u'(x"04"),
u'(x"df"),u'(x"cc"),u'(x"78"),u'(x"00"),u'(x"97"),u'(x"fe"),u'(x"06"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"cd"),u'(x"78"),u'(x"00"),u'(x"d2"),u'(x"b1"),u'(x"02"),
u'(x"04"),u'(x"df"),u'(x"ce"),u'(x"78"),u'(x"00"),u'(x"17"),u'(x"04"),u'(x"04"),u'(x"df"),u'(x"cf"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"0a"),u'(x"57"),u'(x"9c"),
u'(x"cb"),u'(x"77"),u'(x"96"),u'(x"ff"),u'(x"ff"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"fa"),u'(x"00"),u'(x"09"),u'(x"00"),u'(x"03"),u'(x"ff"),u'(x"ff"),u'(x"08"),
u'(x"01"),u'(x"ff"),u'(x"ff"),u'(x"2e"),u'(x"01"),u'(x"d2"),u'(x"96"),u'(x"88"),u'(x"00"),u'(x"04"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"a9"),u'(x"04"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"04"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"08"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"01"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"08"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"00"),u'(x"2a"),u'(x"57"),u'(x"01"),u'(x"46"),u'(x"b5"),u'(x"07"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"02"),
u'(x"00"),u'(x"09"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"ff"),u'(x"09"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"ff"),u'(x"08"),u'(x"ff"),u'(x"ff"),u'(x"1f"),u'(x"fe"),
u'(x"06"),u'(x"c5"),u'(x"00"),u'(x"c1"),u'(x"02"),u'(x"df"),u'(x"5f"),u'(x"00"),u'(x"df"),u'(x"c8"),u'(x"02"),u'(x"bf"),u'(x"97"),u'(x"02"),u'(x"c6"),u'(x"fe"),
u'(x"df"),u'(x"d0"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"06"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"d1"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"bc"),
u'(x"84"),u'(x"06"),u'(x"06"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"d2"),u'(x"78"),u'(x"00"),u'(x"5f"),u'(x"00"),u'(x"5f"),u'(x"02"),u'(x"c6"),u'(x"fe"),u'(x"c2"),
u'(x"06"),u'(x"c3"),u'(x"27"),u'(x"bf"),u'(x"c2"),u'(x"df"),u'(x"02"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"d3"),u'(x"78"),u'(x"00"),u'(x"c2"),u'(x"06"),u'(x"04"),
u'(x"df"),u'(x"d4"),u'(x"78"),u'(x"00"),u'(x"c3"),u'(x"27"),u'(x"04"),u'(x"df"),u'(x"d5"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"c5"),u'(x"04"),u'(x"bf"),u'(x"17"),
u'(x"00"),u'(x"df"),u'(x"07"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"d6"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"d7"),u'(x"78"),u'(x"00"),
u'(x"c5"),u'(x"04"),u'(x"04"),u'(x"df"),u'(x"d8"),u'(x"78"),u'(x"00"),u'(x"c0"),u'(x"04"),u'(x"c5"),u'(x"08"),u'(x"04"),u'(x"bf"),u'(x"00"),u'(x"df"),u'(x"00"),
u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"d9"),u'(x"78"),u'(x"00"),u'(x"c0"),u'(x"04"),u'(x"04"),u'(x"df"),u'(x"da"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"02"),u'(x"04"),
u'(x"df"),u'(x"db"),u'(x"78"),u'(x"00"),u'(x"c5"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"dc"),u'(x"78"),u'(x"00"),u'(x"c5"),u'(x"08"),u'(x"04"),u'(x"bf"),u'(x"17"),
u'(x"03"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"dd"),u'(x"78"),u'(x"00"),u'(x"c4"),u'(x"02"),u'(x"04"),u'(x"df"),u'(x"de"),u'(x"78"),u'(x"00"),
u'(x"c5"),u'(x"02"),u'(x"04"),u'(x"df"),u'(x"df"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"64"),u'(x"5f"),u'(x"ca"),u'(x"44"),u'(x"43"),u'(x"04"),u'(x"45"),u'(x"02"),
u'(x"bf"),u'(x"31"),u'(x"04"),u'(x"5f"),u'(x"06"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"e0"),u'(x"78"),u'(x"00"),u'(x"45"),u'(x"08"),u'(x"04"),u'(x"df"),u'(x"e1"),
u'(x"78"),u'(x"00"),u'(x"44"),u'(x"0a"),u'(x"04"),u'(x"df"),u'(x"e2"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"ca"),u'(x"06"),u'(x"df"),u'(x"e3"),u'(x"78"),u'(x"00"),
u'(x"c1"),u'(x"ca"),u'(x"43"),u'(x"04"),u'(x"06"),u'(x"df"),u'(x"e4"),u'(x"78"),u'(x"00"),u'(x"f1"),u'(x"04"),u'(x"c1"),u'(x"0c"),u'(x"57"),u'(x"db"),u'(x"c9"),
u'(x"77"),u'(x"ce"),u'(x"ff"),u'(x"ff"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"0a"),u'(x"ff"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"ff"),u'(x"02"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"a2"),u'(x"a3"),u'(x"04"),u'(x"a2"),u'(x"00"),u'(x"00"),u'(x"5f"),u'(x"63"),u'(x"04"),u'(x"5f"),u'(x"00"),
u'(x"00"),u'(x"a3"),u'(x"a3"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"fe"),u'(x"11"),u'(x"0a"),u'(x"fe"),u'(x"00"),u'(x"c0"),u'(x"1b"),u'(x"11"),u'(x"08"),
u'(x"c7"),u'(x"14"),u'(x"c0"),u'(x"1b"),u'(x"ef"),u'(x"00"),u'(x"c7"),u'(x"ec"),u'(x"00"),u'(x"ff"),u'(x"01"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"ff"),u'(x"ce"),
u'(x"01"),u'(x"0a"),u'(x"ce"),u'(x"ff"),u'(x"00"),u'(x"02"),u'(x"f8"),u'(x"04"),u'(x"02"),u'(x"00"),u'(x"ff"),u'(x"fe"),u'(x"08"),u'(x"04"),u'(x"fe"),u'(x"00"),
u'(x"01"),u'(x"ff"),u'(x"01"),u'(x"02"),u'(x"ff"),u'(x"01"),u'(x"01"),u'(x"00"),u'(x"02"),u'(x"02"),u'(x"00"),u'(x"01"),u'(x"01"),u'(x"00"),u'(x"03"),u'(x"00"),
u'(x"01"),u'(x"55"),u'(x"13"),u'(x"2c"),u'(x"5f"),u'(x"00"),u'(x"92"),u'(x"a6"),u'(x"db"),u'(x"1f"),u'(x"fe"),u'(x"c2"),u'(x"01"),u'(x"bf"),u'(x"82"),u'(x"df"),
u'(x"00"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"e5"),u'(x"78"),u'(x"00"),u'(x"97"),u'(x"02"),u'(x"04"),u'(x"df"),u'(x"e6"),u'(x"78"),u'(x"00"),u'(x"c2"),u'(x"00"),
u'(x"c3"),u'(x"01"),u'(x"af"),u'(x"83"),u'(x"df"),u'(x"07"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"e7"),u'(x"78"),u'(x"00"),u'(x"d7"),u'(x"01"),u'(x"04"),u'(x"df"),
u'(x"e8"),u'(x"78"),u'(x"00"),u'(x"97"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"e9"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"e6"),u'(x"43"),u'(x"42"),u'(x"02"),u'(x"bf"),
u'(x"89"),u'(x"5f"),u'(x"04"),u'(x"fe"),u'(x"04"),u'(x"df"),u'(x"ea"),u'(x"78"),u'(x"00"),u'(x"42"),u'(x"06"),u'(x"04"),u'(x"df"),u'(x"eb"),u'(x"78"),u'(x"00"),
u'(x"c1"),u'(x"04"),u'(x"df"),u'(x"ec"),u'(x"78"),u'(x"00"),u'(x"c9"),u'(x"04"),u'(x"df"),u'(x"ed"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"08"),u'(x"57"),u'(x"86"),
u'(x"db"),u'(x"77"),u'(x"a0"),u'(x"f1"),u'(x"ff"),u'(x"05"),u'(x"00"),u'(x"c0"),u'(x"ff"),u'(x"00"),u'(x"ff"),u'(x"c0"),u'(x"00"),u'(x"08"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"08"),u'(x"00"),u'(x"df"),u'(x"ff"),u'(x"09"),u'(x"ff"),u'(x"c6"),u'(x"00"),u'(x"07"),u'(x"00"),u'(x"c8"),u'(x"ff"),u'(x"0b"),u'(x"00"),u'(x"cb"),
u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"c7"),u'(x"01"),u'(x"02"),u'(x"80"),u'(x"cf"),u'(x"01"),u'(x"0a"),u'(x"00"),u'(x"e0"),u'(x"ff"),u'(x"04"),u'(x"00"),u'(x"f9"),
u'(x"00"),u'(x"08"),u'(x"a0"),u'(x"e2"),u'(x"00"),u'(x"09"),u'(x"ff"),u'(x"f4"),u'(x"00"),u'(x"08"),u'(x"f8"),u'(x"e8"),u'(x"55"),u'(x"04"),u'(x"00"),u'(x"f0"),
u'(x"00"),u'(x"09"),u'(x"ff"),u'(x"f8"),u'(x"00"),u'(x"08"),u'(x"80"),u'(x"ca"),u'(x"f7"),u'(x"0b"),u'(x"00"),u'(x"f4"),u'(x"ff"),u'(x"01"),u'(x"01"),u'(x"c1"),
u'(x"00"),u'(x"03"),u'(x"00"),u'(x"1f"),u'(x"fe"),u'(x"c1"),u'(x"13"),u'(x"c5"),u'(x"55"),u'(x"04"),u'(x"bf"),u'(x"01"),u'(x"d7"),u'(x"fe"),u'(x"0a"),u'(x"04"),
u'(x"df"),u'(x"ee"),u'(x"78"),u'(x"00"),u'(x"57"),u'(x"13"),u'(x"04"),u'(x"df"),u'(x"ef"),u'(x"78"),u'(x"00"),u'(x"17"),u'(x"a8"),u'(x"04"),u'(x"df"),u'(x"f0"),
u'(x"78"),u'(x"00"),u'(x"57"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"f1"),u'(x"78"),u'(x"00"),u'(x"c3"),u'(x"55"),u'(x"02"),u'(x"c4"),u'(x"d9"),u'(x"bf"),u'(x"d7"),
u'(x"13"),u'(x"d7"),u'(x"fe"),u'(x"0a"),u'(x"04"),u'(x"df"),u'(x"f2"),u'(x"78"),u'(x"00"),u'(x"97"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"f3"),u'(x"78"),u'(x"00"),
u'(x"d7"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"f4"),u'(x"78"),u'(x"00"),u'(x"17"),u'(x"d9"),u'(x"04"),u'(x"df"),u'(x"f5"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"80"),
u'(x"44"),u'(x"42"),u'(x"02"),u'(x"43"),u'(x"04"),u'(x"bf"),u'(x"89"),u'(x"f1"),u'(x"fe"),u'(x"06"),u'(x"04"),u'(x"df"),u'(x"f6"),u'(x"78"),u'(x"00"),u'(x"42"),
u'(x"08"),u'(x"04"),u'(x"df"),u'(x"f7"),u'(x"78"),u'(x"00"),u'(x"43"),u'(x"0a"),u'(x"04"),u'(x"df"),u'(x"f8"),u'(x"78"),u'(x"00"),u'(x"01"),u'(x"04"),u'(x"df"),
u'(x"f9"),u'(x"78"),u'(x"00"),u'(x"4c"),u'(x"04"),u'(x"df"),u'(x"fa"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"0c"),u'(x"57"),u'(x"88"),u'(x"d2"),u'(x"77"),u'(x"08"),
u'(x"c0"),u'(x"55"),u'(x"ff"),u'(x"08"),u'(x"55"),u'(x"ff"),u'(x"ff"),u'(x"01"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"c1"),u'(x"ff"),u'(x"00"),u'(x"0a"),
u'(x"ff"),u'(x"00"),u'(x"c6"),u'(x"ae"),u'(x"c0"),u'(x"02"),u'(x"bf"),u'(x"00"),u'(x"c9"),u'(x"c0"),u'(x"0a"),u'(x"0b"),u'(x"00"),u'(x"00"),u'(x"df"),u'(x"00"),
u'(x"01"),u'(x"04"),u'(x"00"),u'(x"00"),u'(x"de"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"e0"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"ff"),u'(x"ff"),
u'(x"d5"),u'(x"ff"),u'(x"00"),u'(x"07"),u'(x"00"),u'(x"00"),u'(x"d4"),u'(x"ff"),u'(x"00"),u'(x"09"),u'(x"00"),u'(x"00"),u'(x"db"),u'(x"ff"),u'(x"13"),u'(x"0a"),
u'(x"00"),u'(x"00"),u'(x"d7"),u'(x"00"),u'(x"ff"),u'(x"0b"),u'(x"80"),u'(x"00"),u'(x"cf"),u'(x"ff"),u'(x"01"),u'(x"09"),u'(x"00"),u'(x"00"),u'(x"e1"),u'(x"00"),
u'(x"00"),u'(x"08"),u'(x"ff"),u'(x"ff"),u'(x"e2"),u'(x"ff"),u'(x"ff"),u'(x"05"),u'(x"00"),u'(x"00"),u'(x"e2"),u'(x"ff"),u'(x"ff"),u'(x"01"),u'(x"00"),u'(x"01"),
u'(x"c9"),u'(x"80"),u'(x"0a"),u'(x"03"),u'(x"00"),u'(x"00"),u'(x"e0"),u'(x"ff"),u'(x"ff"),u'(x"04"),u'(x"00"),u'(x"00"),u'(x"df"),u'(x"ff"),u'(x"fc"),u'(x"09"),
u'(x"ff"),u'(x"ff"),u'(x"e7"),u'(x"00"),u'(x"00"),u'(x"08"),u'(x"ff"),u'(x"c0"),u'(x"eb"),u'(x"d4"),u'(x"02"),u'(x"01"),u'(x"00"),u'(x"66"),u'(x"f5"),u'(x"e9"),
u'(x"99"),u'(x"09"),u'(x"f0"),u'(x"3f"),u'(x"06"),u'(x"b7"),u'(x"3c"),u'(x"c6"),u'(x"02"),u'(x"04"),u'(x"df"),u'(x"fb"),u'(x"78"),u'(x"00"),u'(x"06"),u'(x"b7"),
u'(x"28"),u'(x"b7"),u'(x"24"),u'(x"c6"),u'(x"04"),u'(x"04"),u'(x"df"),u'(x"fc"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"fe"),u'(x"b7"),u'(x"0e"),u'(x"c6"),u'(x"fc"),
u'(x"04"),u'(x"df"),u'(x"fd"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"fe"),u'(x"b7"),u'(x"f8"),u'(x"b7"),u'(x"f4"),u'(x"c6"),u'(x"fa"),u'(x"04"),u'(x"df"),u'(x"fe"),
u'(x"78"),u'(x"00"),u'(x"06"),u'(x"d6"),u'(x"97"),u'(x"02"),u'(x"04"),u'(x"df"),u'(x"ff"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"fe"),u'(x"e6"),u'(x"c6"),u'(x"fc"),
u'(x"04"),u'(x"df"),u'(x"00"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"fe"),u'(x"1f"),u'(x"f6"),u'(x"c6"),u'(x"68"),u'(x"f7"),u'(x"04"),u'(x"a8"),u'(x"df"),u'(x"40"),
u'(x"04"),u'(x"c1"),u'(x"66"),u'(x"c2"),u'(x"64"),u'(x"c3"),u'(x"62"),u'(x"1f"),u'(x"66"),u'(x"26"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"01"),u'(x"78"),u'(x"00"),
u'(x"df"),u'(x"08"),u'(x"f6"),u'(x"03"),u'(x"97"),u'(x"62"),u'(x"04"),u'(x"df"),u'(x"02"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"f6"),u'(x"df"),u'(x"66"),u'(x"04"),
u'(x"5f"),u'(x"66"),u'(x"9f"),u'(x"64"),u'(x"df"),u'(x"62"),u'(x"c6"),u'(x"fe"),u'(x"1f"),u'(x"f6"),u'(x"c6"),u'(x"00"),u'(x"f7"),u'(x"04"),u'(x"46"),u'(x"df"),
u'(x"96"),u'(x"04"),u'(x"1f"),u'(x"fe"),u'(x"26"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"03"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"f6"),u'(x"c5"),u'(x"00"),u'(x"c6"),
u'(x"00"),u'(x"df"),u'(x"b6"),u'(x"04"),u'(x"a5"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"04"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"f6"),u'(x"c6"),u'(x"68"),u'(x"df"),
u'(x"d2"),u'(x"04"),u'(x"66"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"05"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"f6"),u'(x"df"),u'(x"ea"),u'(x"04"),u'(x"c6"),u'(x"fe"),
u'(x"1f"),u'(x"f6"),u'(x"c6"),u'(x"00"),u'(x"f7"),u'(x"08"),u'(x"d6"),u'(x"df"),u'(x"04"),u'(x"08"),u'(x"f7"),u'(x"04"),u'(x"cc"),u'(x"df"),u'(x"10"),u'(x"04"),
u'(x"3f"),u'(x"a0"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"06"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"b2"),u'(x"04"),u'(x"df"),u'(x"aa"),u'(x"08"),u'(x"1f"),u'(x"f6"),
u'(x"c6"),u'(x"fe"),u'(x"1f"),u'(x"f6"),u'(x"c6"),u'(x"00"),u'(x"f7"),u'(x"10"),u'(x"92"),u'(x"df"),u'(x"48"),u'(x"10"),u'(x"f7"),u'(x"04"),u'(x"88"),u'(x"df"),
u'(x"54"),u'(x"04"),u'(x"04"),u'(x"a0"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"07"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"f6"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"66"),
u'(x"04"),u'(x"df"),u'(x"5e"),u'(x"10"),u'(x"1f"),u'(x"f6"),u'(x"c6"),u'(x"00"),u'(x"f7"),u'(x"18"),u'(x"4e"),u'(x"df"),u'(x"8c"),u'(x"18"),u'(x"f7"),u'(x"04"),
u'(x"44"),u'(x"df"),u'(x"98"),u'(x"04"),u'(x"00"),u'(x"a0"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"08"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"28"),u'(x"18"),u'(x"df"),
u'(x"24"),u'(x"04"),u'(x"1f"),u'(x"f6"),u'(x"c6"),u'(x"fe"),u'(x"1f"),u'(x"f6"),u'(x"c6"),u'(x"00"),u'(x"f7"),u'(x"1c"),u'(x"0a"),u'(x"df"),u'(x"d0"),u'(x"1c"),
u'(x"f7"),u'(x"04"),u'(x"00"),u'(x"df"),u'(x"dc"),u'(x"04"),u'(x"00"),u'(x"a0"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"09"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"e4"),
u'(x"1c"),u'(x"df"),u'(x"e0"),u'(x"04"),u'(x"1f"),u'(x"f6"),u'(x"c6"),u'(x"fe"),u'(x"1f"),u'(x"f6"),u'(x"c6"),u'(x"00"),u'(x"f7"),u'(x"0c"),u'(x"c6"),u'(x"df"),
u'(x"14"),u'(x"0c"),u'(x"f7"),u'(x"04"),u'(x"bc"),u'(x"df"),u'(x"20"),u'(x"04"),u'(x"03"),u'(x"a0"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"0a"),u'(x"78"),u'(x"00"),
u'(x"1f"),u'(x"f6"),u'(x"df"),u'(x"9c"),u'(x"0c"),u'(x"df"),u'(x"98"),u'(x"04"),u'(x"c6"),u'(x"fe"),u'(x"1f"),u'(x"f6"),u'(x"c6"),u'(x"00"),u'(x"f7"),u'(x"08"),
u'(x"82"),u'(x"df"),u'(x"5a"),u'(x"08"),u'(x"f7"),u'(x"04"),u'(x"78"),u'(x"df"),u'(x"66"),u'(x"04"),u'(x"01"),u'(x"41"),u'(x"a0"),u'(x"c6"),u'(x"fe"),u'(x"df"),
u'(x"0b"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"5c"),u'(x"04"),u'(x"df"),u'(x"54"),u'(x"08"),u'(x"1f"),u'(x"f6"),u'(x"c6"),u'(x"fe"),u'(x"1f"),u'(x"f6"),u'(x"c6"),
u'(x"00"),u'(x"f7"),u'(x"08"),u'(x"3c"),u'(x"df"),u'(x"9a"),u'(x"08"),u'(x"df"),u'(x"a6"),u'(x"04"),u'(x"01"),u'(x"41"),u'(x"a0"),u'(x"c6"),u'(x"fe"),u'(x"df"),
u'(x"0c"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"f6"),u'(x"df"),u'(x"16"),u'(x"08"),u'(x"df"),u'(x"12"),u'(x"04"),u'(x"c6"),u'(x"fe"),u'(x"f7"),u'(x"04"),u'(x"04"),
u'(x"df"),u'(x"e0"),u'(x"04"),u'(x"c6"),u'(x"02"),u'(x"e6"),u'(x"c6"),u'(x"02"),u'(x"e6"),u'(x"c6"),u'(x"02"),u'(x"e6"),u'(x"c6"),u'(x"02"),u'(x"e6"),u'(x"06"),
u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"0d"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"d4"),u'(x"04"),u'(x"c6"),u'(x"fe"),u'(x"c6"),u'(x"fe"),u'(x"f7"),u'(x"0c"),u'(x"c4"),
u'(x"e6"),u'(x"10"),u'(x"e6"),u'(x"18"),u'(x"df"),u'(x"20"),u'(x"0c"),u'(x"02"),u'(x"df"),u'(x"0e"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"0f"),u'(x"78"),u'(x"00"),
u'(x"c6"),u'(x"fa"),u'(x"04"),u'(x"df"),u'(x"10"),u'(x"78"),u'(x"00"),u'(x"97"),u'(x"18"),u'(x"04"),u'(x"df"),u'(x"11"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"84"),
u'(x"0c"),u'(x"c6"),u'(x"fe"),u'(x"c6"),u'(x"fe"),u'(x"f7"),u'(x"0c"),u'(x"74"),u'(x"e6"),u'(x"10"),u'(x"e6"),u'(x"68"),u'(x"df"),u'(x"72"),u'(x"0c"),u'(x"06"),
u'(x"df"),u'(x"12"),u'(x"78"),u'(x"00"),u'(x"a0"),u'(x"df"),u'(x"13"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"fa"),u'(x"04"),u'(x"df"),u'(x"14"),u'(x"78"),u'(x"00"),
u'(x"97"),u'(x"6a"),u'(x"04"),u'(x"df"),u'(x"15"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"32"),u'(x"0c"),u'(x"c6"),u'(x"fe"),u'(x"c6"),u'(x"fe"),u'(x"f7"),u'(x"0c"),
u'(x"22"),u'(x"e6"),u'(x"10"),u'(x"e6"),u'(x"c2"),u'(x"df"),u'(x"ca"),u'(x"0c"),u'(x"df"),u'(x"ef"),u'(x"fe"),u'(x"bf"),u'(x"02"),u'(x"df"),u'(x"16"),u'(x"78"),
u'(x"00"),u'(x"df"),u'(x"17"),u'(x"78"),u'(x"00"),u'(x"d7"),u'(x"2e"),u'(x"10"),u'(x"04"),u'(x"df"),u'(x"18"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"fe"),u'(x"e6"),
u'(x"ff"),u'(x"e6"),u'(x"fe"),u'(x"df"),u'(x"06"),u'(x"0c"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"af"),u'(x"02"),u'(x"df"),u'(x"19"),u'(x"78"),u'(x"00"),u'(x"df"),
u'(x"1a"),u'(x"78"),u'(x"00"),u'(x"d7"),u'(x"f2"),u'(x"ff"),u'(x"04"),u'(x"df"),u'(x"1b"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"aa"),u'(x"0c"),u'(x"c6"),u'(x"fe"),
u'(x"c6"),u'(x"fe"),u'(x"f7"),u'(x"08"),u'(x"9a"),u'(x"df"),u'(x"3a"),u'(x"08"),u'(x"3f"),u'(x"df"),u'(x"1c"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"fa"),u'(x"04"),
u'(x"df"),u'(x"1d"),u'(x"78"),u'(x"00"),u'(x"97"),u'(x"32"),u'(x"04"),u'(x"df"),u'(x"1e"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"6a"),u'(x"08"),u'(x"c6"),u'(x"fe"),
u'(x"c6"),u'(x"fe"),u'(x"f7"),u'(x"08"),u'(x"5a"),u'(x"df"),u'(x"80"),u'(x"08"),u'(x"1f"),u'(x"fe"),u'(x"af"),u'(x"3f"),u'(x"df"),u'(x"1f"),u'(x"78"),u'(x"00"),
u'(x"d7"),u'(x"78"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"20"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"ac"),u'(x"08"),u'(x"df"),u'(x"ef"),u'(x"fe"),
u'(x"bf"),u'(x"3f"),u'(x"df"),u'(x"21"),u'(x"78"),u'(x"00"),u'(x"d7"),u'(x"4c"),u'(x"ef"),u'(x"04"),u'(x"df"),u'(x"22"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"04"),
u'(x"08"),u'(x"c6"),u'(x"fe"),u'(x"c6"),u'(x"fe"),u'(x"f7"),u'(x"1c"),u'(x"f4"),u'(x"df"),u'(x"e6"),u'(x"1c"),u'(x"1f"),u'(x"fe"),u'(x"af"),u'(x"00"),u'(x"df"),
u'(x"23"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"fa"),u'(x"04"),u'(x"df"),u'(x"24"),u'(x"78"),u'(x"00"),u'(x"97"),u'(x"de"),u'(x"04"),u'(x"df"),u'(x"25"),u'(x"78"),
u'(x"00"),u'(x"df"),u'(x"be"),u'(x"1c"),u'(x"c6"),u'(x"fe"),u'(x"c6"),u'(x"fe"),u'(x"f7"),u'(x"1c"),u'(x"ae"),u'(x"df"),u'(x"2c"),u'(x"1c"),u'(x"1f"),u'(x"fe"),
u'(x"af"),u'(x"00"),u'(x"df"),u'(x"26"),u'(x"78"),u'(x"00"),u'(x"d7"),u'(x"cc"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"27"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"fe"),
u'(x"df"),u'(x"58"),u'(x"1c"),u'(x"df"),u'(x"ef"),u'(x"fe"),u'(x"bf"),u'(x"00"),u'(x"df"),u'(x"28"),u'(x"78"),u'(x"00"),u'(x"d7"),u'(x"a0"),u'(x"ef"),u'(x"04"),
u'(x"df"),u'(x"29"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"58"),u'(x"1c"),u'(x"c6"),u'(x"fe"),u'(x"03"),u'(x"c6"),u'(x"fe"),u'(x"f7"),u'(x"1c"),u'(x"46"),u'(x"f7"),
u'(x"04"),u'(x"42"),u'(x"df"),u'(x"a2"),u'(x"04"),u'(x"df"),u'(x"aa"),u'(x"1c"),u'(x"77"),u'(x"16"),u'(x"00"),u'(x"df"),u'(x"2a"),u'(x"78"),u'(x"00"),u'(x"77"),
u'(x"08"),u'(x"df"),u'(x"2b"),u'(x"78"),u'(x"00"),u'(x"83"),u'(x"c6"),u'(x"fe"),u'(x"d7"),u'(x"00"),u'(x"06"),u'(x"df"),u'(x"00"),u'(x"94"),u'(x"df"),u'(x"94"),
u'(x"e9"),u'(x"df"),u'(x"fe"),u'(x"1c"),u'(x"df"),u'(x"fa"),u'(x"04"),u'(x"c6"),u'(x"fe"),u'(x"c6"),u'(x"fe"),u'(x"f7"),u'(x"10"),u'(x"e8"),u'(x"df"),u'(x"ec"),
u'(x"10"),u'(x"04"),u'(x"df"),u'(x"2c"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"fa"),u'(x"04"),u'(x"df"),u'(x"2d"),u'(x"78"),u'(x"00"),u'(x"97"),u'(x"e4"),u'(x"04"),
u'(x"df"),u'(x"2e"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"b8"),u'(x"10"),u'(x"c6"),u'(x"fe"),u'(x"c6"),u'(x"fe"),u'(x"f7"),u'(x"10"),u'(x"a8"),u'(x"df"),u'(x"32"),
u'(x"10"),u'(x"1f"),u'(x"fe"),u'(x"af"),u'(x"04"),u'(x"df"),u'(x"2f"),u'(x"78"),u'(x"00"),u'(x"d7"),u'(x"c6"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"30"),u'(x"78"),
u'(x"00"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"5e"),u'(x"10"),u'(x"df"),u'(x"ef"),u'(x"fe"),u'(x"bf"),u'(x"04"),u'(x"df"),u'(x"31"),u'(x"78"),u'(x"00"),u'(x"d7"),
u'(x"9a"),u'(x"ef"),u'(x"04"),u'(x"df"),u'(x"32"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"52"),u'(x"10"),u'(x"c6"),u'(x"fe"),u'(x"c6"),u'(x"fe"),u'(x"f7"),u'(x"18"),
u'(x"42"),u'(x"df"),u'(x"92"),u'(x"18"),u'(x"00"),u'(x"df"),u'(x"33"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"fa"),u'(x"04"),u'(x"df"),u'(x"34"),u'(x"78"),u'(x"00"),
u'(x"97"),u'(x"8a"),u'(x"04"),u'(x"df"),u'(x"35"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"12"),u'(x"18"),u'(x"c6"),u'(x"fe"),u'(x"c6"),u'(x"fe"),u'(x"f7"),u'(x"18"),
u'(x"02"),u'(x"df"),u'(x"d8"),u'(x"18"),u'(x"1f"),u'(x"fe"),u'(x"af"),u'(x"00"),u'(x"df"),u'(x"36"),u'(x"78"),u'(x"00"),u'(x"d7"),u'(x"20"),u'(x"00"),u'(x"04"),
u'(x"df"),u'(x"37"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"04"),u'(x"18"),u'(x"df"),u'(x"ef"),u'(x"fe"),u'(x"bf"),u'(x"00"),u'(x"df"),u'(x"38"),
u'(x"78"),u'(x"00"),u'(x"d7"),u'(x"f4"),u'(x"ef"),u'(x"04"),u'(x"df"),u'(x"39"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"ac"),u'(x"18"),u'(x"c6"),u'(x"fe"),u'(x"c6"),
u'(x"fe"),u'(x"f7"),u'(x"0c"),u'(x"9c"),u'(x"df"),u'(x"38"),u'(x"0c"),u'(x"03"),u'(x"df"),u'(x"3a"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"fa"),u'(x"04"),u'(x"df"),
u'(x"3b"),u'(x"78"),u'(x"00"),u'(x"97"),u'(x"30"),u'(x"04"),u'(x"df"),u'(x"3c"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"6c"),u'(x"0c"),u'(x"c6"),u'(x"fe"),u'(x"c6"),
u'(x"fe"),u'(x"f7"),u'(x"0c"),u'(x"5c"),u'(x"df"),u'(x"7e"),u'(x"0c"),u'(x"1f"),u'(x"fe"),u'(x"af"),u'(x"03"),u'(x"df"),u'(x"3d"),u'(x"78"),u'(x"00"),u'(x"d7"),
u'(x"7a"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"3e"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"aa"),u'(x"0c"),u'(x"df"),u'(x"ef"),u'(x"fe"),u'(x"bf"),
u'(x"03"),u'(x"df"),u'(x"3f"),u'(x"78"),u'(x"00"),u'(x"d7"),u'(x"4e"),u'(x"ef"),u'(x"04"),u'(x"df"),u'(x"40"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"06"),u'(x"0c"),
u'(x"c6"),u'(x"fe"),u'(x"c6"),u'(x"fe"),u'(x"f7"),u'(x"08"),u'(x"f6"),u'(x"df"),u'(x"e0"),u'(x"08"),u'(x"01"),u'(x"41"),u'(x"df"),u'(x"41"),u'(x"78"),u'(x"00"),
u'(x"c6"),u'(x"fa"),u'(x"04"),u'(x"df"),u'(x"42"),u'(x"78"),u'(x"00"),u'(x"97"),u'(x"d8"),u'(x"04"),u'(x"df"),u'(x"43"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"c4"),
u'(x"08"),u'(x"c6"),u'(x"fe"),u'(x"c6"),u'(x"fe"),u'(x"f7"),u'(x"08"),u'(x"b4"),u'(x"df"),u'(x"28"),u'(x"08"),u'(x"1f"),u'(x"fe"),u'(x"af"),u'(x"01"),u'(x"41"),
u'(x"df"),u'(x"44"),u'(x"78"),u'(x"00"),u'(x"d7"),u'(x"d0"),u'(x"04"),u'(x"04"),u'(x"df"),u'(x"45"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"54"),
u'(x"08"),u'(x"df"),u'(x"ef"),u'(x"fe"),u'(x"bf"),u'(x"41"),u'(x"df"),u'(x"46"),u'(x"78"),u'(x"00"),u'(x"d7"),u'(x"a4"),u'(x"ef"),u'(x"04"),u'(x"df"),u'(x"47"),
u'(x"78"),u'(x"00"),u'(x"df"),u'(x"5c"),u'(x"08"),u'(x"c6"),u'(x"fe"),u'(x"c6"),u'(x"fe"),u'(x"f7"),u'(x"08"),u'(x"4c"),u'(x"df"),u'(x"8a"),u'(x"08"),u'(x"03"),
u'(x"c3"),u'(x"df"),u'(x"48"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"fa"),u'(x"04"),u'(x"df"),u'(x"49"),u'(x"78"),u'(x"00"),u'(x"97"),u'(x"82"),u'(x"04"),u'(x"df"),
u'(x"4a"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"1a"),u'(x"08"),u'(x"c6"),u'(x"fe"),u'(x"c6"),u'(x"fe"),u'(x"f7"),u'(x"08"),u'(x"0a"),u'(x"df"),u'(x"d2"),u'(x"08"),
u'(x"1f"),u'(x"fe"),u'(x"af"),u'(x"03"),u'(x"c3"),u'(x"df"),u'(x"4b"),u'(x"78"),u'(x"00"),u'(x"d7"),u'(x"26"),u'(x"04"),u'(x"04"),u'(x"df"),u'(x"4c"),u'(x"78"),
u'(x"00"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"fe"),u'(x"08"),u'(x"df"),u'(x"ef"),u'(x"fe"),u'(x"bf"),u'(x"c3"),u'(x"df"),u'(x"4d"),u'(x"78"),u'(x"00"),u'(x"d7"),
u'(x"fa"),u'(x"ef"),u'(x"04"),u'(x"df"),u'(x"4e"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"b2"),u'(x"08"),u'(x"c6"),u'(x"fe"),u'(x"1f"),u'(x"f6"),u'(x"f7"),u'(x"04"),
u'(x"a2"),u'(x"df"),u'(x"3a"),u'(x"04"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"df"),u'(x"c0"),u'(x"df"),u'(x"4f"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"10"),u'(x"f6"),
u'(x"04"),u'(x"df"),u'(x"50"),u'(x"78"),u'(x"00"),u'(x"97"),u'(x"32"),u'(x"04"),u'(x"df"),u'(x"51"),u'(x"78"),u'(x"00"),u'(x"97"),u'(x"00"),u'(x"04"),u'(x"df"),
u'(x"52"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"f6"),u'(x"df"),u'(x"56"),u'(x"04"),u'(x"1f"),u'(x"f6"),u'(x"f7"),u'(x"04"),u'(x"4a"),u'(x"df"),u'(x"9c"),u'(x"04"),
u'(x"f7"),u'(x"06"),u'(x"40"),u'(x"1f"),u'(x"06"),u'(x"e6"),u'(x"00"),u'(x"e6"),u'(x"95"),u'(x"02"),u'(x"df"),u'(x"53"),u'(x"78"),u'(x"00"),u'(x"df"),u'(x"40"),
u'(x"f6"),u'(x"04"),u'(x"df"),u'(x"54"),u'(x"78"),u'(x"00"),u'(x"d6"),u'(x"95"),u'(x"04"),u'(x"df"),u'(x"55"),u'(x"78"),u'(x"00"),u'(x"d6"),u'(x"00"),u'(x"04"),
u'(x"df"),u'(x"56"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"f6"),u'(x"df"),u'(x"e8"),u'(x"04"),u'(x"df"),u'(x"e0"),u'(x"06"),u'(x"1f"),u'(x"fe"),u'(x"5f"),u'(x"fe"),
u'(x"df"),u'(x"57"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"fe"),u'(x"df"),u'(x"40"),u'(x"f6"),u'(x"04"),u'(x"df"),u'(x"58"),u'(x"78"),u'(x"00"),u'(x"d6"),u'(x"fe"),
u'(x"04"),u'(x"df"),u'(x"59"),u'(x"78"),u'(x"00"),u'(x"d6"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"5a"),u'(x"78"),u'(x"00"),u'(x"c1"),u'(x"e0"),u'(x"04"),u'(x"df"),
u'(x"5b"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"f6"),u'(x"df"),u'(x"96"),u'(x"04"),u'(x"df"),u'(x"92"),u'(x"06"),u'(x"f7"),u'(x"04"),u'(x"88"),u'(x"df"),u'(x"5a"),
u'(x"04"),u'(x"c6"),u'(x"ff"),u'(x"1f"),u'(x"f6"),u'(x"1f"),u'(x"fe"),u'(x"df"),u'(x"c0"),u'(x"df"),u'(x"5c"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"00"),u'(x"04"),
u'(x"df"),u'(x"5d"),u'(x"78"),u'(x"00"),u'(x"d6"),u'(x"52"),u'(x"04"),u'(x"df"),u'(x"5e"),u'(x"78"),u'(x"00"),u'(x"ce"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"5f"),
u'(x"78"),u'(x"00"),u'(x"df"),u'(x"54"),u'(x"f6"),u'(x"04"),u'(x"df"),u'(x"60"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"f6"),u'(x"c6"),u'(x"fe"),u'(x"df"),u'(x"24"),
u'(x"04"),u'(x"1f"),u'(x"00"),u'(x"1f"),u'(x"02"),u'(x"f7"),u'(x"04"),u'(x"14"),u'(x"df"),u'(x"c6"),u'(x"04"),u'(x"1f"),u'(x"f6"),u'(x"df"),u'(x"fa"),u'(x"df"),
u'(x"02"),u'(x"04"),u'(x"04"),u'(x"df"),u'(x"61"),u'(x"78"),u'(x"00"),u'(x"f7"),u'(x"a0"),u'(x"f0"),u'(x"f7"),u'(x"a2"),u'(x"ec"),u'(x"df"),u'(x"88"),u'(x"a0"),
u'(x"df"),u'(x"e0"),u'(x"a2"),u'(x"c3"),u'(x"00"),u'(x"c4"),u'(x"1a"),u'(x"9f"),u'(x"1f"),u'(x"fa"),u'(x"d4"),u'(x"fa"),u'(x"04"),u'(x"df"),u'(x"62"),u'(x"78"),
u'(x"00"),u'(x"df"),u'(x"fa"),u'(x"d4"),u'(x"fa"),u'(x"04"),u'(x"df"),u'(x"63"),u'(x"78"),u'(x"00"),u'(x"c3"),u'(x"f5"),u'(x"08"),u'(x"00"),u'(x"22"),u'(x"44"),
u'(x"66"),u'(x"88"),u'(x"aa"),u'(x"cc"),u'(x"ee"),u'(x"9f"),u'(x"1f"),u'(x"fa"),u'(x"c3"),u'(x"00"),u'(x"c4"),u'(x"56"),u'(x"df"),u'(x"fa"),u'(x"cc"),u'(x"fa"),
u'(x"04"),u'(x"df"),u'(x"64"),u'(x"78"),u'(x"00"),u'(x"03"),u'(x"c3"),u'(x"ff"),u'(x"d4"),u'(x"f2"),u'(x"0c"),u'(x"ee"),u'(x"cc"),u'(x"aa"),u'(x"88"),u'(x"66"),
u'(x"44"),u'(x"22"),u'(x"00"),u'(x"df"),u'(x"65"),u'(x"78"),u'(x"00"),u'(x"c3"),u'(x"00"),u'(x"df"),u'(x"9a"),u'(x"a0"),u'(x"df"),u'(x"e0"),u'(x"a2"),u'(x"04"),
u'(x"d4"),u'(x"df"),u'(x"fa"),u'(x"98"),u'(x"df"),u'(x"66"),u'(x"78"),u'(x"00"),u'(x"c6"),u'(x"04"),u'(x"c3"),u'(x"f4"),u'(x"0e"),u'(x"c5"),u'(x"fa"),u'(x"1f"),
u'(x"fa"),u'(x"c5"),u'(x"f1"),u'(x"05"),u'(x"04"),u'(x"df"),u'(x"67"),u'(x"78"),u'(x"00"),u'(x"77"),u'(x"da"),u'(x"1f"),u'(x"fa"),u'(x"1f"),u'(x"fe"),u'(x"9f"),
u'(x"c3"),u'(x"00"),u'(x"df"),u'(x"de"),u'(x"a0"),u'(x"df"),u'(x"e0"),u'(x"a2"),u'(x"df"),u'(x"fa"),u'(x"c3"),u'(x"fc"),u'(x"1f"),u'(x"fa"),u'(x"06"),u'(x"1f"),
u'(x"fa"),u'(x"df"),u'(x"68"),u'(x"78"),u'(x"00"),u'(x"1f"),u'(x"fa"),u'(x"df"),u'(x"3e"),u'(x"a0"),u'(x"df"),u'(x"e0"),u'(x"a2"),u'(x"c5"),u'(x"78"),u'(x"df") 
);
signal memo : mem_type := mem_type'(
u'(x"00"),u'(x"01"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"15"),u'(x"01"),u'(x"00"),u'(x"2b"),u'(x"0a"),u'(x"53"),u'(x"17"),u'(x"53"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"03"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"02"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"86"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),
u'(x"87"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"02"),u'(x"0a"),u'(x"02"),u'(x"0b"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"15"),u'(x"aa"),u'(x"00"),u'(x"25"),u'(x"aa"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),u'(x"00"),u'(x"27"),u'(x"00"),
u'(x"55"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"27"),u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"ff"),u'(x"20"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"20"),u'(x"00"),u'(x"03"),u'(x"15"),
u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"20"),u'(x"aa"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),u'(x"20"),u'(x"55"),
u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"ff"),u'(x"20"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"20"),
u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"20"),u'(x"aa"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),
u'(x"55"),u'(x"20"),u'(x"55"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"ff"),u'(x"20"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"0a"),u'(x"20"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"20"),u'(x"aa"),u'(x"03"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),u'(x"20"),u'(x"55"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"ff"),u'(x"20"),u'(x"ff"),u'(x"03"),
u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"20"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"20"),u'(x"aa"),
u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),u'(x"20"),u'(x"55"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"ff"),
u'(x"21"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"21"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),
u'(x"aa"),u'(x"21"),u'(x"aa"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),u'(x"21"),u'(x"55"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"15"),u'(x"ff"),u'(x"21"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"21"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"21"),u'(x"aa"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),u'(x"21"),u'(x"55"),u'(x"03"),
u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"ff"),u'(x"21"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"21"),u'(x"00"),
u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"21"),u'(x"aa"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),
u'(x"21"),u'(x"55"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"25"),u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"25"),u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"25"),
u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"25"),u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"8a"),u'(x"80"),u'(x"8a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"03"),u'(x"80"),u'(x"0a"),u'(x"03"),u'(x"15"),
u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"8a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"8a"),u'(x"81"),u'(x"03"),
u'(x"8a"),u'(x"8a"),u'(x"8a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"03"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"8a"),u'(x"80"),u'(x"03"),u'(x"8a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),
u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"80"),u'(x"0a"),u'(x"0a"),
u'(x"0a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"0a"),u'(x"8a"),u'(x"80"),u'(x"0a"),u'(x"8a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),
u'(x"0a"),u'(x"8a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"8a"),u'(x"80"),u'(x"0a"),u'(x"8a"),u'(x"03"),u'(x"15"),
u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"0a"),
u'(x"80"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),
u'(x"8a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"8a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),
u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"02"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"03"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"8a"),u'(x"0a"),
u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"03"),u'(x"81"),u'(x"0a"),u'(x"0a"),
u'(x"0a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),
u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"8a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"03"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"03"),u'(x"0a"),u'(x"8a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),
u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0b"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"0a"),u'(x"0b"),u'(x"03"),u'(x"85"),u'(x"81"),u'(x"87"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"8a"),u'(x"0b"),u'(x"03"),u'(x"85"),u'(x"86"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"8a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"00"),u'(x"03"),u'(x"15"),
u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"01"),u'(x"03"),u'(x"0a"),u'(x"01"),u'(x"0a"),u'(x"01"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),
u'(x"0a"),u'(x"0b"),u'(x"00"),u'(x"03"),u'(x"85"),u'(x"81"),u'(x"87"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"0b"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"8b"),u'(x"00"),u'(x"85"),u'(x"03"),u'(x"80"),u'(x"87"),u'(x"15"),
u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"8a"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),
u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),
u'(x"00"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"01"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),
u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"0b"),u'(x"ff"),u'(x"87"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0b"),u'(x"01"),u'(x"03"),
u'(x"85"),u'(x"81"),u'(x"87"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"0b"),u'(x"87"),u'(x"85"),u'(x"81"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"00"),
u'(x"0b"),u'(x"87"),u'(x"85"),u'(x"03"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"8a"),u'(x"00"),u'(x"00"),u'(x"8b"),u'(x"85"),u'(x"87"),
u'(x"85"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"8b"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"00"),
u'(x"00"),u'(x"0b"),u'(x"87"),u'(x"85"),u'(x"81"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0b"),u'(x"03"),u'(x"85"),u'(x"87"),
u'(x"80"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"8b"),u'(x"87"),u'(x"85"),u'(x"81"),u'(x"03"),
u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"8b"),u'(x"03"),u'(x"81"),u'(x"85"),u'(x"86"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),
u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"0b"),u'(x"87"),u'(x"85"),u'(x"81"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0b"),
u'(x"87"),u'(x"85"),u'(x"03"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"8b"),u'(x"85"),
u'(x"87"),u'(x"81"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"8b"),u'(x"03"),u'(x"87"),u'(x"85"),u'(x"81"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"0b"),u'(x"87"),u'(x"85"),u'(x"81"),u'(x"03"),u'(x"15"),
u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"0b"),u'(x"87"),u'(x"03"),u'(x"85"),u'(x"81"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"00"),u'(x"0b"),u'(x"87"),u'(x"85"),u'(x"81"),u'(x"03"),
u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"0b"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),
u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"8b"),u'(x"03"),u'(x"87"),u'(x"85"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"0a"),u'(x"0a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"0b"),u'(x"87"),u'(x"85"),
u'(x"81"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0b"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),
u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8b"),u'(x"03"),u'(x"87"),u'(x"85"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"8b"),u'(x"03"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"0b"),u'(x"87"),u'(x"85"),u'(x"81"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0b"),
u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"8b"),u'(x"87"),u'(x"81"),u'(x"85"),
u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"8b"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),
u'(x"0a"),u'(x"0a"),u'(x"0b"),u'(x"ff"),u'(x"87"),u'(x"85"),u'(x"81"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0b"),u'(x"01"),u'(x"03"),
u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"0a"),u'(x"0b"),u'(x"ff"),
u'(x"87"),u'(x"85"),u'(x"03"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0b"),u'(x"ff"),u'(x"81"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"10"),u'(x"03"),u'(x"85"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"02"),u'(x"0a"),u'(x"0a"),
u'(x"0a"),u'(x"60"),u'(x"03"),u'(x"87"),u'(x"85"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"e0"),u'(x"85"),u'(x"86"),u'(x"03"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"e0"),u'(x"03"),
u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"03"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),u'(x"81"),
u'(x"02"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"60"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"02"),u'(x"0a"),u'(x"0a"),u'(x"15"),
u'(x"aa"),u'(x"15"),u'(x"55"),u'(x"00"),u'(x"40"),u'(x"86"),u'(x"85"),u'(x"03"),u'(x"80"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"21"),u'(x"03"),u'(x"15"),
u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"50"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"02"),u'(x"15"),u'(x"aa"),
u'(x"15"),u'(x"80"),u'(x"15"),u'(x"55"),u'(x"31"),u'(x"03"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"21"),u'(x"03"),u'(x"86"),u'(x"81"),u'(x"15"),
u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"20"),u'(x"03"),u'(x"87"),u'(x"85"),u'(x"80"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"00"),u'(x"31"),
u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"8a"),u'(x"0a"),u'(x"15"),u'(x"01"),
u'(x"00"),u'(x"13"),u'(x"03"),u'(x"85"),u'(x"86"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"02"),u'(x"00"),u'(x"92"),u'(x"03"),u'(x"81"),
u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"8a"),u'(x"02"),u'(x"0a"),u'(x"92"),u'(x"80"),u'(x"85"),u'(x"87"),u'(x"25"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"ff"),u'(x"15"),u'(x"00"),u'(x"62"),u'(x"03"),u'(x"87"),u'(x"80"),u'(x"0a"),u'(x"03"),
u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"e3"),u'(x"03"),u'(x"81"),
u'(x"86"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"e3"),u'(x"02"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"55"),u'(x"15"),u'(x"aa"),u'(x"53"),
u'(x"03"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"43"),u'(x"03"),u'(x"81"),
u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"42"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"55"),u'(x"15"),
u'(x"01"),u'(x"15"),u'(x"aa"),u'(x"00"),u'(x"33"),u'(x"87"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"23"),u'(x"03"),u'(x"86"),u'(x"84"),u'(x"81"),
u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"32"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),
u'(x"15"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0b"),u'(x"00"),u'(x"14"),u'(x"81"),u'(x"86"),u'(x"85"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"0a"),u'(x"63"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"ff"),u'(x"15"),u'(x"ff"),u'(x"e5"),
u'(x"03"),u'(x"85"),u'(x"86"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"e5"),u'(x"ff"),u'(x"81"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"c3"),u'(x"15"),u'(x"ff"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"ff"),u'(x"45"),
u'(x"03"),u'(x"80"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"55"),u'(x"c5"),u'(x"0a"),u'(x"d5"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),
u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"aa"),u'(x"15"),u'(x"80"),u'(x"15"),u'(x"80"),u'(x"0b"),
u'(x"b5"),u'(x"81"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"b4"),u'(x"03"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"03"),
u'(x"86"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0b"),u'(x"24"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"15"),
u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"58"),u'(x"ef"),u'(x"00"),u'(x"03"),u'(x"87"),u'(x"80"),
u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"58"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"15"),
u'(x"aa"),u'(x"15"),u'(x"f6"),u'(x"29"),u'(x"87"),u'(x"80"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"00"),u'(x"b8"),u'(x"86"),u'(x"03"),
u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0b"),u'(x"0a"),u'(x"a9"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"00"),
u'(x"15"),u'(x"ff"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"6b"),u'(x"03"),u'(x"80"),u'(x"86"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"65"),u'(x"00"),u'(x"6a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"aa"),u'(x"15"),u'(x"00"),u'(x"15"),
u'(x"80"),u'(x"3d"),u'(x"01"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"bd"),u'(x"01"),u'(x"ff"),u'(x"03"),u'(x"81"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"0a"),u'(x"15"),u'(x"ff"),u'(x"15"),u'(x"ff"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"0a"),u'(x"ef"),u'(x"fe"),
u'(x"01"),u'(x"03"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"ee"),u'(x"ff"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),
u'(x"aa"),u'(x"00"),u'(x"0c"),u'(x"84"),u'(x"86"),u'(x"25"),u'(x"55"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"00"),u'(x"8c"),
u'(x"86"),u'(x"84"),u'(x"81"),u'(x"25"),u'(x"aa"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"15"),u'(x"55"),u'(x"0c"),u'(x"80"),u'(x"84"),
u'(x"87"),u'(x"23"),u'(x"aa"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"0a"),u'(x"00"),u'(x"8c"),u'(x"81"),u'(x"86"),u'(x"84"),
u'(x"0a"),u'(x"25"),u'(x"55"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"15"),u'(x"80"),u'(x"00"),u'(x"0c"),u'(x"86"),u'(x"84"),u'(x"03"),
u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"02"),u'(x"15"),u'(x"08"),u'(x"00"),u'(x"8c"),u'(x"87"),u'(x"85"),u'(x"0a"),u'(x"25"),u'(x"08"),
u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"15"),u'(x"55"),u'(x"00"),u'(x"0c"),u'(x"00"),u'(x"80"),u'(x"84"),u'(x"87"),u'(x"25"),u'(x"aa"),
u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"00"),u'(x"8c"),u'(x"00"),u'(x"81"),u'(x"86"),u'(x"85"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"0a"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"58"),u'(x"00"),u'(x"0c"),u'(x"80"),u'(x"84"),u'(x"87"),u'(x"25"),u'(x"b1"),u'(x"02"),u'(x"0b"),u'(x"03"),
u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"a7"),u'(x"00"),u'(x"0c"),u'(x"81"),u'(x"86"),u'(x"84"),u'(x"0b"),u'(x"02"),
u'(x"25"),u'(x"4e"),u'(x"01"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"0a"),u'(x"15"),u'(x"35"),u'(x"00"),u'(x"0c"),u'(x"ff"),
u'(x"81"),u'(x"87"),u'(x"85"),u'(x"25"),u'(x"6a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"0a"),u'(x"01"),u'(x"15"),u'(x"80"),
u'(x"00"),u'(x"0c"),u'(x"00"),u'(x"81"),u'(x"02"),u'(x"86"),u'(x"84"),u'(x"0b"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),
u'(x"15"),u'(x"41"),u'(x"00"),u'(x"01"),u'(x"81"),u'(x"25"),u'(x"c0"),u'(x"02"),u'(x"00"),u'(x"01"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),
u'(x"55"),u'(x"00"),u'(x"0c"),u'(x"86"),u'(x"25"),u'(x"2a"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"8c"),
u'(x"86"),u'(x"80"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"52"),u'(x"15"),u'(x"12"),u'(x"00"),u'(x"27"),
u'(x"52"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"20"),u'(x"12"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"52"),
u'(x"15"),u'(x"12"),u'(x"00"),u'(x"12"),u'(x"27"),u'(x"52"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"52"),u'(x"15"),u'(x"12"),
u'(x"00"),u'(x"27"),u'(x"52"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"12"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"0a"),u'(x"52"),u'(x"15"),u'(x"12"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"13"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"27"),u'(x"52"),u'(x"00"),
u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"52"),u'(x"15"),u'(x"12"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"12"),u'(x"03"),u'(x"15"),
u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"27"),u'(x"52"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"52"),u'(x"15"),u'(x"13"),u'(x"00"),
u'(x"12"),u'(x"25"),u'(x"00"),u'(x"52"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"52"),u'(x"15"),u'(x"13"),u'(x"00"),u'(x"ff"),u'(x"13"),
u'(x"00"),u'(x"25"),u'(x"00"),u'(x"52"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"13"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),
u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),
u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),
u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),
u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),
u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),
u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"14"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"13"),u'(x"15"),u'(x"00"),u'(x"65"),u'(x"00"),u'(x"7e"),u'(x"15"),u'(x"00"),u'(x"52"),u'(x"00"),u'(x"0b"),u'(x"52"),
u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"52"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"27"),u'(x"52"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"52"),u'(x"00"),u'(x"14"),u'(x"27"),u'(x"52"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"52"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"14"),u'(x"27"),u'(x"52"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"27"),u'(x"52"),u'(x"00"),
u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"52"),u'(x"00"),u'(x"ff"),u'(x"15"),u'(x"01"),u'(x"11"),u'(x"52"),u'(x"11"),u'(x"52"),u'(x"e5"),
u'(x"00"),u'(x"52"),u'(x"15"),u'(x"00"),u'(x"52"),u'(x"15"),u'(x"14"),u'(x"0a"),u'(x"0a"),u'(x"09"),u'(x"25"),u'(x"00"),u'(x"52"),u'(x"03"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"27"),u'(x"52"),u'(x"02"),u'(x"23"),u'(x"aa"),u'(x"02"),u'(x"25"),u'(x"15"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),
u'(x"52"),u'(x"17"),u'(x"52"),u'(x"15"),u'(x"14"),u'(x"0a"),u'(x"09"),u'(x"00"),u'(x"15"),u'(x"25"),u'(x"00"),u'(x"52"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"27"),u'(x"52"),u'(x"02"),u'(x"23"),u'(x"ff"),u'(x"02"),u'(x"25"),u'(x"14"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"52"),
u'(x"17"),u'(x"52"),u'(x"15"),u'(x"aa"),u'(x"15"),u'(x"14"),u'(x"09"),u'(x"25"),u'(x"00"),u'(x"52"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"27"),
u'(x"52"),u'(x"02"),u'(x"23"),u'(x"55"),u'(x"02"),u'(x"25"),u'(x"15"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"52"),u'(x"17"),u'(x"52"),
u'(x"15"),u'(x"00"),u'(x"15"),u'(x"15"),u'(x"09"),u'(x"00"),u'(x"15"),u'(x"25"),u'(x"00"),u'(x"52"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"27"),
u'(x"52"),u'(x"02"),u'(x"23"),u'(x"00"),u'(x"02"),u'(x"25"),u'(x"14"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"52"),u'(x"17"),u'(x"52"),
u'(x"15"),u'(x"55"),u'(x"15"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"25"),u'(x"00"),u'(x"52"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"27"),u'(x"52"),
u'(x"02"),u'(x"23"),u'(x"a7"),u'(x"02"),u'(x"25"),u'(x"16"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"52"),u'(x"17"),u'(x"52"),u'(x"15"),
u'(x"ff"),u'(x"15"),u'(x"15"),u'(x"09"),u'(x"ff"),u'(x"16"),u'(x"25"),u'(x"00"),u'(x"52"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"27"),u'(x"52"),
u'(x"02"),u'(x"23"),u'(x"00"),u'(x"02"),u'(x"25"),u'(x"15"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"52"),u'(x"17"),u'(x"52"),u'(x"15"),
u'(x"a7"),u'(x"15"),u'(x"15"),u'(x"09"),u'(x"ff"),u'(x"25"),u'(x"00"),u'(x"52"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"27"),u'(x"52"),u'(x"02"),
u'(x"23"),u'(x"ff"),u'(x"02"),u'(x"25"),u'(x"15"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"17"),u'(x"52"),u'(x"15"),u'(x"00"),u'(x"52"),u'(x"11"),
u'(x"52"),u'(x"11"),u'(x"52"),u'(x"e5"),u'(x"00"),u'(x"52"),u'(x"15"),u'(x"ff"),u'(x"09"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"52"),u'(x"02"),u'(x"27"),u'(x"52"),
u'(x"02"),u'(x"23"),u'(x"ff"),u'(x"02"),u'(x"21"),u'(x"16"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"52"),u'(x"15"),u'(x"d5"),u'(x"17"),
u'(x"52"),u'(x"09"),u'(x"16"),u'(x"00"),u'(x"27"),u'(x"52"),u'(x"00"),u'(x"02"),u'(x"27"),u'(x"52"),u'(x"02"),u'(x"23"),u'(x"00"),u'(x"02"),u'(x"21"),u'(x"17"),
u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"52"),u'(x"17"),u'(x"52"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"00"),u'(x"00"),u'(x"17"),u'(x"27"),
u'(x"52"),u'(x"00"),u'(x"02"),u'(x"27"),u'(x"52"),u'(x"02"),u'(x"23"),u'(x"d5"),u'(x"02"),u'(x"21"),u'(x"16"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"0a"),u'(x"52"),u'(x"17"),u'(x"52"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"ff"),u'(x"27"),u'(x"52"),u'(x"00"),u'(x"02"),u'(x"27"),u'(x"52"),u'(x"02"),u'(x"23"),
u'(x"00"),u'(x"02"),u'(x"21"),u'(x"16"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"17"),u'(x"52"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"a7"),u'(x"15"),
u'(x"17"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"a7"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"11"),u'(x"15"),u'(x"17"),
u'(x"11"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"23"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"10"),u'(x"15"),u'(x"40"),u'(x"ff"),
u'(x"15"),u'(x"ff"),u'(x"25"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"25"),u'(x"aa"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),u'(x"25"),u'(x"55"),u'(x"03"),u'(x"15"),
u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"c0"),u'(x"ff"),u'(x"15"),u'(x"ff"),u'(x"25"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"0a"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"25"),u'(x"aa"),u'(x"03"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),u'(x"25"),u'(x"55"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"0a"),u'(x"ff"),u'(x"15"),
u'(x"01"),u'(x"0a"),u'(x"01"),u'(x"0a"),u'(x"01"),u'(x"0a"),u'(x"01"),u'(x"09"),u'(x"00"),u'(x"15"),u'(x"40"),u'(x"ff"),u'(x"25"),u'(x"01"),u'(x"03"),u'(x"15"),
u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"c0"),u'(x"ff"),u'(x"25"),u'(x"01"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"25"),
u'(x"01"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"40"),u'(x"ff"),u'(x"09"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),
u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"c0"),u'(x"ff"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),
u'(x"25"),u'(x"18"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"c0"),u'(x"ff"),u'(x"09"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),
u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"25"),u'(x"18"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"40"),u'(x"ff"),
u'(x"25"),u'(x"18"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"18"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),
u'(x"40"),u'(x"ff"),u'(x"25"),u'(x"18"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"25"),u'(x"18"),u'(x"03"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"c0"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"81"),u'(x"85"),u'(x"86"),u'(x"03"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"80"),u'(x"03"),u'(x"85"),u'(x"87"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),
u'(x"00"),u'(x"00"),u'(x"35"),u'(x"00"),u'(x"81"),u'(x"85"),u'(x"86"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"35"),u'(x"80"),
u'(x"03"),u'(x"85"),u'(x"87"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"45"),u'(x"ff"),u'(x"81"),u'(x"85"),
u'(x"86"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"45"),u'(x"7f"),u'(x"03"),u'(x"85"),u'(x"87"),u'(x"81"),u'(x"15"),
u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"55"),u'(x"00"),u'(x"81"),u'(x"85"),u'(x"86"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"55"),u'(x"80"),u'(x"03"),u'(x"85"),u'(x"87"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"7f"),u'(x"00"),u'(x"00"),
u'(x"0a"),u'(x"03"),u'(x"80"),u'(x"84"),u'(x"87"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"0a"),u'(x"87"),u'(x"85"),u'(x"0a"),u'(x"85"),u'(x"87"),
u'(x"00"),u'(x"00"),u'(x"0a"),u'(x"03"),u'(x"84"),u'(x"86"),u'(x"80"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"0a"),u'(x"81"),u'(x"85"),
u'(x"87"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0b"),u'(x"03"),u'(x"85"),u'(x"87"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"85"),u'(x"87"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"7f"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"61"),
u'(x"84"),u'(x"87"),u'(x"03"),u'(x"81"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"61"),u'(x"84"),u'(x"86"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"61"),u'(x"85"),u'(x"87"),u'(x"81"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"ff"),u'(x"00"),u'(x"0b"),u'(x"81"),u'(x"85"),u'(x"86"),
u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"7f"),u'(x"00"),u'(x"00"),u'(x"0b"),u'(x"80"),u'(x"87"),u'(x"03"),u'(x"85"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"0b"),u'(x"85"),u'(x"87"),u'(x"81"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"7f"),u'(x"00"),u'(x"0b"),u'(x"85"),
u'(x"86"),u'(x"03"),u'(x"81"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0b"),u'(x"81"),u'(x"87"),u'(x"85"),u'(x"03"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"7f"),u'(x"15"),u'(x"f0"),u'(x"00"),u'(x"21"),u'(x"84"),u'(x"86"),u'(x"03"),u'(x"81"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),
u'(x"00"),u'(x"0a"),u'(x"81"),u'(x"03"),u'(x"86"),u'(x"84"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"0a"),u'(x"81"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"15"),u'(x"7f"),u'(x"00"),u'(x"e5"),u'(x"bf"),u'(x"84"),u'(x"80"),u'(x"03"),u'(x"87"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"00"),
u'(x"00"),u'(x"e5"),u'(x"00"),u'(x"86"),u'(x"85"),u'(x"03"),u'(x"81"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"80"),u'(x"00"),u'(x"0b"),u'(x"80"),
u'(x"85"),u'(x"00"),u'(x"0b"),u'(x"84"),u'(x"87"),u'(x"80"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"0b"),u'(x"87"),u'(x"85"),
u'(x"02"),u'(x"00"),u'(x"0b"),u'(x"86"),u'(x"85"),u'(x"03"),u'(x"81"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"60"),u'(x"00"),u'(x"0c"),u'(x"87"),
u'(x"84"),u'(x"81"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0c"),u'(x"86"),u'(x"85"),u'(x"81"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0c"),u'(x"84"),
u'(x"86"),u'(x"81"),u'(x"02"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0c"),u'(x"85"),u'(x"87"),u'(x"80"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),
u'(x"00"),u'(x"00"),u'(x"0c"),u'(x"86"),u'(x"84"),u'(x"80"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0c"),u'(x"86"),u'(x"85"),u'(x"81"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"0c"),u'(x"84"),u'(x"87"),u'(x"81"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0c"),u'(x"85"),u'(x"87"),u'(x"80"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),u'(x"00"),u'(x"0c"),u'(x"0c"),u'(x"0c"),u'(x"87"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"4a"),u'(x"03"),
u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"00"),u'(x"0c"),u'(x"0c"),u'(x"0c"),u'(x"87"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),
u'(x"55"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"60"),u'(x"00"),u'(x"0c"),u'(x"87"),u'(x"84"),u'(x"81"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"0c"),u'(x"86"),u'(x"85"),u'(x"81"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0c"),u'(x"84"),u'(x"86"),u'(x"81"),u'(x"03"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"0c"),u'(x"85"),u'(x"87"),u'(x"80"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"0c"),u'(x"86"),u'(x"84"),
u'(x"80"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"55"),u'(x"80"),u'(x"0c"),u'(x"86"),u'(x"85"),u'(x"81"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0c"),
u'(x"84"),u'(x"87"),u'(x"81"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0c"),u'(x"84"),u'(x"87"),u'(x"80"),u'(x"25"),u'(x"f0"),u'(x"03"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"a7"),u'(x"11"),u'(x"00"),u'(x"0d"),u'(x"87"),u'(x"81"),u'(x"85"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"10"),
u'(x"00"),u'(x"0d"),u'(x"03"),u'(x"80"),u'(x"86"),u'(x"85"),u'(x"0a"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"a7"),u'(x"15"),u'(x"55"),
u'(x"00"),u'(x"78"),u'(x"85"),u'(x"03"),u'(x"87"),u'(x"81"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"00"),u'(x"78"),u'(x"81"),u'(x"03"),
u'(x"86"),u'(x"84"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"79"),u'(x"85"),u'(x"81"),u'(x"86"),u'(x"02"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"0d"),u'(x"85"),u'(x"80"),u'(x"03"),u'(x"86"),u'(x"0a"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"0a"),u'(x"15"),u'(x"00"),u'(x"0d"),u'(x"02"),u'(x"85"),u'(x"87"),u'(x"81"),u'(x"0b"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),
u'(x"15"),u'(x"ff"),u'(x"0a"),u'(x"0d"),u'(x"0b"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"15"),u'(x"ff"),u'(x"0d"),u'(x"25"),u'(x"ff"),
u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"0f"),u'(x"15"),u'(x"b6"),u'(x"00"),u'(x"79"),u'(x"80"),u'(x"03"),u'(x"86"),u'(x"85"),u'(x"20"),
u'(x"b9"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"10"),u'(x"00"),u'(x"79"),u'(x"81"),u'(x"85"),u'(x"87"),u'(x"20"),u'(x"0f"),u'(x"03"),u'(x"15"),
u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"00"),u'(x"86"),u'(x"84"),u'(x"80"),u'(x"02"),u'(x"7f"),u'(x"86"),u'(x"84"),u'(x"80"),u'(x"02"),u'(x"00"),
u'(x"00"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"21"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"aa"),u'(x"01"),u'(x"15"),u'(x"1e"),u'(x"15"),u'(x"0d"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"82"),u'(x"80"),u'(x"85"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"aa"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"21"),
u'(x"01"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),u'(x"15"),u'(x"0d"),u'(x"11"),u'(x"09"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"83"),u'(x"81"),u'(x"84"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"21"),u'(x"01"),u'(x"03"),u'(x"15"),
u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"55"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"30"),
u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"30"),
u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"30"),
u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"30"),
u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"30"),
u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),
u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),
u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),
u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),
u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),
u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),
u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),
u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),
u'(x"04"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"06"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"07"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),
u'(x"05"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"07"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"06"),u'(x"01"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"05"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"07"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"04"),u'(x"01"),
u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"06"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"07"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"05"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"04"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"06"),u'(x"01"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"04"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"06"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"07"),u'(x"01"),
u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"05"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"ff"),u'(x"15"),u'(x"00"),u'(x"15"),
u'(x"00"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"11"),u'(x"52"),u'(x"15"),u'(x"30"),u'(x"52"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"09"),u'(x"00"),u'(x"21"),u'(x"52"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"52"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"09"),u'(x"00"),u'(x"21"),u'(x"52"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"27"),u'(x"52"),u'(x"ff"),
u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),
u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),
u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"15"),u'(x"08"),u'(x"ff"),u'(x"35"),u'(x"08"),u'(x"ff"),u'(x"02"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"15"),u'(x"ff"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"11"),u'(x"45"),u'(x"08"),u'(x"ff"),u'(x"35"),u'(x"08"),u'(x"ff"),u'(x"03"),u'(x"15"),
u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0b"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0b"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0b"),
u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0b"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0b"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"0b"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"08"),u'(x"ff"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),
u'(x"45"),u'(x"08"),u'(x"ff"),u'(x"15"),u'(x"ff"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"11"),u'(x"55"),u'(x"08"),u'(x"ff"),u'(x"0b"),u'(x"03"),u'(x"15"),
u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0b"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0b"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0b"),
u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0b"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0b"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"15"),u'(x"ff"),u'(x"20"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"20"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"20"),u'(x"aa"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),u'(x"20"),u'(x"55"),u'(x"03"),
u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"ff"),u'(x"20"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"20"),u'(x"00"),
u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"20"),u'(x"aa"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),
u'(x"20"),u'(x"55"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"ff"),u'(x"20"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),
u'(x"0a"),u'(x"20"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"20"),u'(x"aa"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"15"),u'(x"55"),u'(x"20"),u'(x"55"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"ff"),u'(x"20"),u'(x"ff"),u'(x"03"),u'(x"15"),
u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"20"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"20"),u'(x"aa"),u'(x"03"),
u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),u'(x"20"),u'(x"55"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"ff"),u'(x"21"),
u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"21"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"aa"),
u'(x"21"),u'(x"aa"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),u'(x"21"),u'(x"55"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),
u'(x"15"),u'(x"ff"),u'(x"21"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"21"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"15"),u'(x"aa"),u'(x"21"),u'(x"aa"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),u'(x"21"),u'(x"55"),u'(x"03"),u'(x"15"),
u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"45"),u'(x"08"),u'(x"ff"),u'(x"0a"),u'(x"15"),u'(x"26"),u'(x"15"),u'(x"26"),u'(x"15"),u'(x"26"),u'(x"14"),u'(x"ff"),u'(x"8d"),
u'(x"27"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"21"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"22"),u'(x"ff"),u'(x"02"),
u'(x"15"),u'(x"26"),u'(x"15"),u'(x"26"),u'(x"15"),u'(x"26"),u'(x"11"),u'(x"12"),u'(x"ff"),u'(x"8d"),u'(x"27"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"21"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"11"),u'(x"15"),u'(x"26"),u'(x"15"),u'(x"26"),u'(x"15"),u'(x"26"),u'(x"0a"),u'(x"52"),
u'(x"15"),u'(x"52"),u'(x"14"),u'(x"ff"),u'(x"8d"),u'(x"27"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"21"),u'(x"52"),u'(x"03"),u'(x"15"),
u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"27"),u'(x"52"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"22"),u'(x"ff"),u'(x"02"),u'(x"00"),u'(x"00"),u'(x"30"),
u'(x"30"),u'(x"30"),u'(x"ff"),u'(x"30"),u'(x"30"),u'(x"30"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"ff"),
u'(x"15"),u'(x"27"),u'(x"15"),u'(x"27"),u'(x"10"),u'(x"09"),u'(x"00"),u'(x"15"),u'(x"c0"),u'(x"ff"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"27"),u'(x"15"),u'(x"27"),
u'(x"10"),u'(x"09"),u'(x"00"),u'(x"15"),u'(x"c0"),u'(x"ff"),u'(x"15"),u'(x"27"),u'(x"15"),u'(x"27"),u'(x"15"),u'(x"27"),u'(x"10"),u'(x"09"),u'(x"00"),u'(x"15"),
u'(x"30"),u'(x"ff"),u'(x"15"),u'(x"27"),u'(x"15"),u'(x"27"),u'(x"15"),u'(x"27"),u'(x"0a"),u'(x"ff"),u'(x"8d"),u'(x"ff"),u'(x"25"),u'(x"00"),u'(x"ff"),u'(x"03"),
u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"14"),u'(x"8d"),u'(x"27"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"24"),
u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"22"),u'(x"ff"),u'(x"02"),u'(x"00"),u'(x"8d"),u'(x"27"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"a5"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"20"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"22"),u'(x"ff"),
u'(x"02"),u'(x"00"),u'(x"00"),u'(x"55"),u'(x"30"),u'(x"30"),u'(x"30"),u'(x"ff"),u'(x"c0"),u'(x"c0"),u'(x"c0"),u'(x"c0"),u'(x"ff"),u'(x"ff"),u'(x"ff"),u'(x"ff"),
u'(x"00"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"15"),u'(x"28"),u'(x"00"),u'(x"15"),u'(x"ff"),u'(x"15"),u'(x"30"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),
u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"20"),u'(x"02"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"ff"),u'(x"00"),u'(x"00"),
u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"20"),u'(x"02"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"0a"),u'(x"ff"),u'(x"17"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"17"),
u'(x"00"),u'(x"17"),u'(x"00"),u'(x"15"),u'(x"28"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"15"),u'(x"28"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"15"),u'(x"c0"),u'(x"ff"),
u'(x"15"),u'(x"01"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"25"),u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"28"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"25"),u'(x"c0"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"00"),
u'(x"15"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"ff"),u'(x"15"),u'(x"e0"),u'(x"ff"),u'(x"15"),u'(x"00"),u'(x"f5"),u'(x"0a"),u'(x"ff"),u'(x"27"),u'(x"ff"),u'(x"00"),
u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"2a"),u'(x"ff"),u'(x"25"),u'(x"2a"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),
u'(x"15"),u'(x"7e"),u'(x"ff"),u'(x"25"),u'(x"7e"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"ff"),
u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"17"),u'(x"ff"),u'(x"45"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),
u'(x"25"),u'(x"00"),u'(x"f5"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),
u'(x"17"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"15"),u'(x"29"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"29"),
u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"c0"),u'(x"ff"),u'(x"15"),u'(x"e0"),u'(x"ff"),u'(x"15"),u'(x"00"),u'(x"f5"),u'(x"15"),u'(x"7e"),u'(x"ff"),
u'(x"00"),u'(x"00"),u'(x"25"),u'(x"c0"),u'(x"ff"),u'(x"03"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"17"),u'(x"ff"),u'(x"45"),u'(x"00"),u'(x"25"),
u'(x"e0"),u'(x"03"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"f5"),u'(x"03"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),
u'(x"25"),u'(x"7e"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"0a"),u'(x"ff"),u'(x"10"),u'(x"00"),u'(x"10"),
u'(x"00"),u'(x"11"),u'(x"00"),u'(x"11"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"2a"),u'(x"15"),u'(x"30"),u'(x"ff"),u'(x"09"),u'(x"00"),u'(x"24"),u'(x"ff"),
u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"7f"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"c0"),u'(x"ff"),u'(x"15"),u'(x"01"),u'(x"09"),u'(x"00"),u'(x"25"),
u'(x"c0"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"7f"),u'(x"00"),u'(x"00"),u'(x"21"),u'(x"00"),u'(x"02"),u'(x"00"),u'(x"00"),u'(x"01"),
u'(x"21"),u'(x"00"),u'(x"02"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"21"),u'(x"00"),u'(x"02"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"21"),u'(x"00"),u'(x"02"),u'(x"00"),
u'(x"00"),u'(x"01"),u'(x"21"),u'(x"00"),u'(x"02"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"21"),u'(x"00"),u'(x"02"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"21"),u'(x"00"),
u'(x"02"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"30"),u'(x"30"),u'(x"30"),u'(x"30"),u'(x"30"),u'(x"30"),u'(x"30"),u'(x"30"),u'(x"0a"),
u'(x"ff"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"2b"),u'(x"14"),u'(x"7e"),u'(x"17"),u'(x"00"),u'(x"15"),u'(x"2b"),u'(x"00"),u'(x"0a"),u'(x"15"),
u'(x"01"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"10"),u'(x"15"),u'(x"30"),u'(x"ff"),u'(x"00"),u'(x"0e"),u'(x"24"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"20"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"21"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),
u'(x"55"),u'(x"00"),u'(x"24"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"22"),u'(x"ff"),u'(x"02"),u'(x"15"),u'(x"2b"),u'(x"00"),
u'(x"0e"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"ef"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"30"),u'(x"30"),u'(x"30"),u'(x"ef"),u'(x"00"),
u'(x"00"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0b"),u'(x"0b"),u'(x"15"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),
u'(x"2c"),u'(x"14"),u'(x"7e"),u'(x"17"),u'(x"00"),u'(x"15"),u'(x"2c"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"10"),u'(x"15"),
u'(x"30"),u'(x"ff"),u'(x"12"),u'(x"20"),u'(x"01"),u'(x"03"),u'(x"02"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"00"),u'(x"0e"),u'(x"24"),u'(x"ff"),u'(x"03"),u'(x"15"),
u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"22"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"20"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),
u'(x"00"),u'(x"24"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"22"),u'(x"ff"),u'(x"02"),u'(x"15"),u'(x"2c"),u'(x"00"),u'(x"0e"),
u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"ef"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"ff"),u'(x"ff"),u'(x"30"),u'(x"30"),u'(x"30"),
u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0b"),u'(x"0b"),u'(x"15"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"2d"),u'(x"10"),u'(x"52"),u'(x"65"),u'(x"00"),
u'(x"52"),u'(x"15"),u'(x"a4"),u'(x"12"),u'(x"00"),u'(x"70"),u'(x"00"),u'(x"2c"),u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"2c"),
u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"2c"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"2c"),u'(x"00"),u'(x"26"),
u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"65"),u'(x"00"),u'(x"20"),u'(x"2d"),u'(x"02"),u'(x"15"),u'(x"2d"),u'(x"10"),u'(x"15"),u'(x"01"),u'(x"15"),
u'(x"00"),u'(x"12"),u'(x"00"),u'(x"71"),u'(x"00"),u'(x"2c"),u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"2c"),u'(x"00"),u'(x"03"),
u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"21"),u'(x"01"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0b"),u'(x"22"),u'(x"00"),
u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"21"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"65"),u'(x"00"),u'(x"20"),u'(x"2d"),
u'(x"02"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"0d"),u'(x"80"),u'(x"00"),u'(x"00"),u'(x"f9"),u'(x"ff"),u'(x"7f"),u'(x"00"),
u'(x"80"),u'(x"ff"),u'(x"7f"),u'(x"01"),u'(x"00"),u'(x"fe"),u'(x"00"),u'(x"f6"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"06"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"80"),u'(x"00"),u'(x"00"),u'(x"80"),u'(x"ff"),u'(x"7f"),u'(x"00"),u'(x"00"),u'(x"7f"),u'(x"00"),
u'(x"00"),u'(x"10"),u'(x"00"),u'(x"80"),u'(x"00"),u'(x"03"),u'(x"39"),u'(x"00"),u'(x"6d"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"07"),u'(x"00"),u'(x"00"),
u'(x"80"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"80"),u'(x"7f"),u'(x"00"),u'(x"80"),u'(x"c0"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"0a"),u'(x"ff"),
u'(x"0a"),u'(x"17"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"2d"),u'(x"00"),u'(x"00"),u'(x"73"),u'(x"00"),u'(x"15"),u'(x"01"),
u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"2d"),
u'(x"0c"),u'(x"21"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"11"),u'(x"00"),u'(x"10"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),
u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"72"),u'(x"25"),u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),
u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"73"),
u'(x"00"),u'(x"25"),u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),
u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"73"),u'(x"25"),u'(x"00"),
u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),
u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"73"),
u'(x"00"),u'(x"25"),u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),
u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"2f"),u'(x"10"),u'(x"52"),u'(x"12"),u'(x"1c"),u'(x"00"),u'(x"1c"),u'(x"00"),
u'(x"00"),u'(x"73"),u'(x"00"),u'(x"2c"),u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"2c"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"2c"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"27"),u'(x"52"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),
u'(x"17"),u'(x"52"),u'(x"2c"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"10"),u'(x"00"),u'(x"65"),u'(x"00"),u'(x"22"),u'(x"00"),u'(x"02"),
u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"0f"),u'(x"0f"),u'(x"00"),u'(x"0f"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"0f"),u'(x"0f"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"80"),u'(x"08"),u'(x"10"),u'(x"00"),u'(x"08"),u'(x"80"),u'(x"ff"),u'(x"f0"),u'(x"10"),u'(x"00"),
u'(x"f2"),u'(x"fc"),u'(x"ff"),u'(x"f0"),u'(x"ef"),u'(x"00"),u'(x"f2"),u'(x"03"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"ff"),u'(x"4b"),
u'(x"00"),u'(x"00"),u'(x"4b"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"55"),u'(x"00"),u'(x"1c"),u'(x"1d"),u'(x"00"),u'(x"10"),u'(x"00"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"74"),u'(x"25"),
u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"20"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"80"),
u'(x"15"),u'(x"00"),u'(x"00"),u'(x"74"),u'(x"25"),u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"20"),u'(x"00"),u'(x"03"),u'(x"15"),
u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"20"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"10"),u'(x"1c"),u'(x"00"),u'(x"00"),
u'(x"74"),u'(x"2c"),u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"2c"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),
u'(x"20"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"22"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"65"),u'(x"00"),u'(x"20"),u'(x"31"),
u'(x"02"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"7f"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"1f"),u'(x"00"),u'(x"1f"),u'(x"ff"),u'(x"80"),u'(x"00"),u'(x"80"),u'(x"ff"),
u'(x"80"),u'(x"00"),u'(x"c0"),u'(x"ff"),u'(x"ff"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"84"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"1f"),u'(x"00"),u'(x"ff"),u'(x"ff"),
u'(x"00"),u'(x"00"),u'(x"50"),u'(x"ff"),u'(x"f0"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"80"),u'(x"ff"),u'(x"1f"),u'(x"00"),u'(x"00"),u'(x"ff"),
u'(x"d0"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"80"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"80"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"55"),u'(x"00"),u'(x"00"),u'(x"ff"),
u'(x"80"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"80"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"08"),u'(x"00"),u'(x"dc"),u'(x"ff"),u'(x"1f"),u'(x"00"),u'(x"00"),u'(x"ff"),
u'(x"90"),u'(x"00"),u'(x"20"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"55"),u'(x"0a"),u'(x"00"),u'(x"77"),u'(x"27"),u'(x"ff"),u'(x"00"),u'(x"03"),
u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"20"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"21"),u'(x"aa"),u'(x"03"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"21"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"55"),u'(x"0a"),u'(x"15"),u'(x"e9"),u'(x"00"),u'(x"76"),
u'(x"00"),u'(x"27"),u'(x"ff"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"20"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),
u'(x"20"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"21"),u'(x"e9"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"32"),
u'(x"10"),u'(x"1c"),u'(x"00"),u'(x"1c"),u'(x"00"),u'(x"00"),u'(x"76"),u'(x"27"),u'(x"ff"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"2c"),
u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"2c"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"21"),u'(x"03"),u'(x"15"),
u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"22"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"65"),u'(x"00"),u'(x"20"),u'(x"33"),u'(x"02"),u'(x"00"),u'(x"01"),
u'(x"ff"),u'(x"80"),u'(x"ff"),u'(x"00"),u'(x"80"),u'(x"ff"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"80"),u'(x"ff"),u'(x"4f"),u'(x"80"),u'(x"00"),
u'(x"9f"),u'(x"00"),u'(x"ff"),u'(x"08"),u'(x"ff"),u'(x"00"),u'(x"2b"),u'(x"f0"),u'(x"ff"),u'(x"6b"),u'(x"00"),u'(x"00"),u'(x"80"),u'(x"14"),u'(x"ff"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"40"),u'(x"00"),u'(x"ff"),u'(x"80"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"ff"),
u'(x"ff"),u'(x"ff"),u'(x"f8"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"f8"),u'(x"00"),u'(x"80"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"de"),u'(x"00"),
u'(x"98"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"80"),u'(x"80"),u'(x"ff"),u'(x"80"),
u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"ff"),u'(x"3f"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"7f"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"ff"),u'(x"6b"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"14"),u'(x"ff"),u'(x"7f"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"ff"),u'(x"00"),
u'(x"ff"),u'(x"ff"),u'(x"ff"),u'(x"80"),u'(x"f8"),u'(x"00"),u'(x"ff"),u'(x"ff"),u'(x"ff"),u'(x"0c"),u'(x"72"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"84"),
u'(x"fe"),u'(x"00"),u'(x"ff"),u'(x"9d"),u'(x"0a"),u'(x"95"),u'(x"1f"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"95"),
u'(x"1f"),u'(x"95"),u'(x"1f"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"99"),u'(x"1f"),u'(x"25"),u'(x"01"),
u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"99"),u'(x"1e"),u'(x"99"),u'(x"1e"),u'(x"25"),u'(x"01"),u'(x"03"),u'(x"15"),u'(x"01"),
u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"8b"),u'(x"21"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"01"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"8b"),u'(x"25"),u'(x"01"),
u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"1e"),u'(x"15"),u'(x"34"),
u'(x"00"),u'(x"17"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),
u'(x"25"),u'(x"00"),u'(x"ff"),u'(x"02"),u'(x"21"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"1d"),u'(x"1e"),u'(x"00"),
u'(x"10"),u'(x"00"),u'(x"10"),u'(x"00"),u'(x"10"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"1e"),u'(x"15"),
u'(x"34"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"02"),u'(x"15"),
u'(x"01"),u'(x"15"),u'(x"34"),u'(x"00"),u'(x"69"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"00"),u'(x"15"),
u'(x"34"),u'(x"00"),u'(x"49"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"1d"),u'(x"1d"),u'(x"00"),u'(x"15"),u'(x"01"),
u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"1d"),u'(x"15"),u'(x"35"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"1d"),u'(x"15"),u'(x"35"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"1d"),u'(x"00"),u'(x"1d"),u'(x"1d"),u'(x"00"),u'(x"0a"),u'(x"ff"),
u'(x"15"),u'(x"01"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"1d"),u'(x"15"),u'(x"35"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"1d"),u'(x"15"),
u'(x"35"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"01"),u'(x"1d"),u'(x"1d"),
u'(x"00"),u'(x"1d"),u'(x"1d"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"1d"),u'(x"15"),u'(x"35"),u'(x"00"),u'(x"17"),u'(x"00"),
u'(x"1d"),u'(x"15"),u'(x"35"),u'(x"00"),u'(x"88"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"1d"),u'(x"00"),u'(x"1d"),
u'(x"1d"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"01"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"1d"),u'(x"15"),u'(x"35"),u'(x"00"),
u'(x"17"),u'(x"00"),u'(x"1d"),u'(x"15"),u'(x"35"),u'(x"00"),u'(x"89"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"1c"),
u'(x"00"),u'(x"1d"),u'(x"1c"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"01"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"1c"),u'(x"15"),
u'(x"36"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"1c"),u'(x"15"),u'(x"36"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),
u'(x"0a"),u'(x"ff"),u'(x"1d"),u'(x"1c"),u'(x"00"),u'(x"1d"),u'(x"1c"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),
u'(x"1c"),u'(x"15"),u'(x"36"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"1c"),u'(x"15"),u'(x"36"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),
u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"1c"),u'(x"00"),u'(x"1d"),u'(x"1c"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"01"),u'(x"0a"),u'(x"ff"),u'(x"15"),
u'(x"01"),u'(x"17"),u'(x"00"),u'(x"1c"),u'(x"15"),u'(x"36"),u'(x"00"),u'(x"15"),u'(x"36"),u'(x"00"),u'(x"0a"),u'(x"09"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),
u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"1d"),u'(x"1c"),u'(x"00"),u'(x"1d"),u'(x"1c"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"1c"),
u'(x"15"),u'(x"36"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"0b"),u'(x"15"),u'(x"04"),u'(x"0b"),u'(x"15"),u'(x"08"),u'(x"0b"),u'(x"15"),u'(x"10"),u'(x"0b"),u'(x"01"),
u'(x"15"),u'(x"01"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"1b"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"1b"),
u'(x"15"),u'(x"00"),u'(x"15"),u'(x"37"),u'(x"15"),u'(x"37"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),
u'(x"25"),u'(x"01"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"23"),u'(x"37"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"1b"),
u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"1b"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"37"),u'(x"15"),u'(x"37"),u'(x"00"),u'(x"00"),
u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"01"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),
u'(x"23"),u'(x"37"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"1b"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),
u'(x"1b"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"37"),u'(x"15"),u'(x"37"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),
u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"2d"),u'(x"ca"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),
u'(x"00"),u'(x"15"),u'(x"37"),u'(x"15"),u'(x"38"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"15"),
u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"2d"),u'(x"c9"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"1a"),u'(x"00"),u'(x"15"),u'(x"01"),
u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"1a"),u'(x"15"),u'(x"38"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"01"),u'(x"03"),
u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"23"),u'(x"38"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"1a"),u'(x"00"),u'(x"15"),u'(x"01"),
u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"1a"),u'(x"15"),u'(x"38"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),
u'(x"2d"),u'(x"c9"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"38"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),
u'(x"00"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"2d"),u'(x"c9"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"1a"),
u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"19"),u'(x"15"),u'(x"38"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"00"),u'(x"89"),u'(x"15"),
u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"01"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"23"),u'(x"38"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),
u'(x"00"),u'(x"1d"),u'(x"19"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"19"),u'(x"15"),u'(x"39"),u'(x"00"),u'(x"0a"),u'(x"ff"),
u'(x"00"),u'(x"89"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"2d"),u'(x"c8"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),
u'(x"15"),u'(x"39"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"89"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"2d"),u'(x"c8"),u'(x"00"),u'(x"03"),
u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"19"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"0a"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"19"),u'(x"17"),
u'(x"00"),u'(x"19"),u'(x"15"),u'(x"39"),u'(x"00"),u'(x"15"),u'(x"39"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"15"),u'(x"01"),u'(x"20"),u'(x"01"),u'(x"03"),u'(x"15"),u'(x"89"),u'(x"39"),u'(x"60"),u'(x"39"),
u'(x"01"),u'(x"1d"),u'(x"18"),u'(x"00"),u'(x"1d"),u'(x"18"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"18"),u'(x"15"),u'(x"39"),
u'(x"00"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"01"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"23"),u'(x"39"),u'(x"03"),
u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"18"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"18"),u'(x"15"),u'(x"3a"),
u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"2d"),u'(x"c7"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),
u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"3a"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"2d"),
u'(x"c7"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"18"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),
u'(x"18"),u'(x"15"),u'(x"3a"),u'(x"00"),u'(x"88"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"01"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),
u'(x"23"),u'(x"3a"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"18"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),
u'(x"18"),u'(x"15"),u'(x"3a"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"00"),u'(x"88"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"2d"),u'(x"c7"),u'(x"00"),u'(x"03"),
u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"3b"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"88"),u'(x"15"),u'(x"02"),
u'(x"ff"),u'(x"00"),u'(x"2d"),u'(x"c6"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"17"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),
u'(x"01"),u'(x"17"),u'(x"00"),u'(x"17"),u'(x"15"),u'(x"3b"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"01"),u'(x"03"),u'(x"15"),
u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"23"),u'(x"3b"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"17"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),
u'(x"01"),u'(x"17"),u'(x"00"),u'(x"17"),u'(x"15"),u'(x"3b"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"2d"),
u'(x"c6"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"3b"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),
u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"2d"),u'(x"c6"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"17"),u'(x"00"),
u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"16"),u'(x"15"),u'(x"3b"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),
u'(x"25"),u'(x"01"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"23"),u'(x"3b"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"16"),
u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"16"),u'(x"15"),u'(x"3c"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"00"),
u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"2d"),u'(x"c5"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"3c"),
u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"2d"),u'(x"c5"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"02"),
u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"16"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"16"),u'(x"15"),u'(x"3c"),u'(x"00"),u'(x"0a"),
u'(x"08"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"01"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"23"),u'(x"3c"),u'(x"03"),u'(x"15"),
u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"16"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"01"),u'(x"17"),u'(x"00"),u'(x"16"),u'(x"15"),u'(x"3c"),u'(x"00"),
u'(x"0a"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"08"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"2d"),u'(x"c5"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),
u'(x"00"),u'(x"15"),u'(x"01"),u'(x"15"),u'(x"3c"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"08"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"2d"),
u'(x"c4"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"1d"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"01"),u'(x"0a"),u'(x"ff"),u'(x"17"),u'(x"00"),
u'(x"15"),u'(x"15"),u'(x"3d"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"ff"),u'(x"0b"),u'(x"ff"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"ff"),
u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"3d"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"03"),u'(x"15"),
u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"1d"),u'(x"15"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"17"),u'(x"00"),u'(x"15"),u'(x"15"),u'(x"3d"),u'(x"00"),
u'(x"17"),u'(x"00"),u'(x"15"),u'(x"0a"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"15"),u'(x"3d"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),
u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"3d"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"30"),u'(x"03"),
u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"3d"),u'(x"00"),u'(x"15"),u'(x"30"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"00"),u'(x"ff"),
u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"17"),u'(x"ff"),u'(x"25"),u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"ff"),
u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),
u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"1d"),u'(x"14"),u'(x"00"),u'(x"1d"),u'(x"14"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"14"),u'(x"15"),u'(x"3e"),
u'(x"00"),u'(x"15"),u'(x"01"),u'(x"0a"),u'(x"ff"),u'(x"0a"),u'(x"ff"),u'(x"0b"),u'(x"ff"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),
u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"3e"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"03"),u'(x"15"),u'(x"02"),
u'(x"ff"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"01"),u'(x"1d"),u'(x"14"),
u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"14"),u'(x"15"),u'(x"3e"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"0b"),u'(x"ff"),u'(x"1d"),
u'(x"14"),u'(x"00"),u'(x"01"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"17"),u'(x"00"),u'(x"13"),u'(x"17"),u'(x"00"),u'(x"13"),u'(x"1d"),u'(x"00"),u'(x"00"),
u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"15"),u'(x"3f"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"27"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),
u'(x"00"),u'(x"10"),u'(x"ff"),u'(x"27"),u'(x"ff"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"0c"),u'(x"86"),u'(x"01"),u'(x"00"),u'(x"02"),u'(x"04"),
u'(x"08"),u'(x"10"),u'(x"20"),u'(x"40"),u'(x"80"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"fe"),u'(x"15"),u'(x"3f"),u'(x"10"),u'(x"ff"),u'(x"27"),u'(x"ff"),
u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"0c"),u'(x"45"),u'(x"01"),u'(x"0b"),u'(x"02"),u'(x"01"),u'(x"fe"),u'(x"7e"),u'(x"3e"),u'(x"1e"),u'(x"0e"),
u'(x"06"),u'(x"02"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"15"),u'(x"3f"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"0a"),
u'(x"0b"),u'(x"50"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"65"),u'(x"00"),u'(x"0c"),u'(x"86"),u'(x"01"),u'(x"17"),u'(x"ff"),u'(x"0a"),
u'(x"ff"),u'(x"45"),u'(x"ff"),u'(x"21"),u'(x"03"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"0a"),u'(x"ff"),u'(x"0a"),u'(x"ff"),u'(x"00"),
u'(x"15"),u'(x"02"),u'(x"15"),u'(x"3f"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"10"),u'(x"ff"),u'(x"0c"),u'(x"86"),u'(x"0a"),u'(x"ff"),u'(x"01"),u'(x"0a"),
u'(x"ff"),u'(x"15"),u'(x"02"),u'(x"ff"),u'(x"00"),u'(x"0a"),u'(x"ff"),u'(x"15"),u'(x"40"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"40"),u'(x"15") 
);


begin
   base_addr_match <= '1' when base_addr(17 downto 14) = bus_addr(17 downto 14) else '0';
   bus_addr_match <= base_addr_match;

   process(clk, base_addr_match)
   begin
      if clk = '1' and clk'event then
         bus_dati(7 downto 0) <= meme(conv_integer(bus_addr(13 downto 1)));
         bus_dati(15 downto 8) <= memo(conv_integer(bus_addr(13 downto 1)));
      end if;
   end process;

   process(clk, base_addr_match)
   begin
      if clk = '1' and clk'event then
         if base_addr_match = '1' and bus_control_dato = '1' then
            if bus_control_datob = '0' or (bus_control_datob = '1' and bus_addr(0) = '0') then
               meme(conv_integer(bus_addr(13 downto 1))) <= bus_dato(7 downto 0);
            end if;
            if bus_control_datob = '0' or (bus_control_datob = '1' and bus_addr(0) = '1') then
               memo(conv_integer(bus_addr(13 downto 1))) <= bus_dato(15 downto 8);
            end if;
         end if;
      end if;
   end process;
end implementation;

